// JPEG Encoder Block
/* Made by D. Krishna Swaroop, 2017A3PS0315P as part of Study oriented Project in 6th Semester
   BITS Pilani. */
  

// This block is the Stimulus Block. TESTBENCH 
`timescale 1ps / 1ps

module jpeg_top_tb;


reg end_of_file_signal;
reg [23:0]data_in;
reg clk;
reg rst;
reg enable;
wire [31:0]JPEG_bitstream;
wire data_ready;
wire [4:0]end_of_file_bitstream_count;
wire eof_data_partial_ready;



// Unit Under Test 
	jpeg_top UUT (
		.end_of_file_signal(end_of_file_signal),
		.data_in(data_in),
		.clk(clk),
		.rst(rst),
		.enable(enable),
		.JPEG_bitstream(JPEG_bitstream),
		.data_ready(data_ready),
		.end_of_file_bitstream_count(end_of_file_bitstream_count),
		.eof_data_partial_ready(eof_data_partial_ready));



initial
begin : STIMUL 
	#0
	rst = 1'b1;
	enable = 1'b0;
	end_of_file_signal = 1'b0;
    #10000; 
	rst = 1'b0;
	enable = 1'b1;
	// data_in holds the red, green, and blue pixel values
	// obtained from the .tif image file. These values will have to changed based o input image. The following are bits values obtained from the Bitmap of the input image.
    
	
	data_in <= 24'b001101100101001101101110;
#10000;
data_in <= 24'b001101110101010001101111;
#10000;
data_in <= 24'b010001110110010001111111;
#10000;
data_in <= 24'b010110100111011110010010;
#10000;
data_in <= 24'b011001011000000010011011;
#10000;
data_in <= 24'b011010001000001110011110;
#10000;
data_in <= 24'b011001000111101110010101;
#10000;
data_in <= 24'b010101100110110010000101;
#10000;
data_in <= 24'b001110010101011001110001;
#10000;
data_in <= 24'b010000000101110101111000;
#10000;
data_in <= 24'b010100010110111010001001;
#10000;
data_in <= 24'b010111000111100110010100;
#10000;
data_in <= 24'b011000000111101110010110;
#10000;
data_in <= 24'b011010011000000110011101;
#10000;
data_in <= 24'b011011101000010110011111;
#10000;
data_in <= 24'b011001110111110110010110;
#10000;
data_in <= 24'b010100110110111010001001;
#10000;
data_in <= 24'b010110100111010110010000;
#10000;
data_in <= 24'b011001000111111110011010;
#10000;
data_in <= 24'b011001000111111110011010;
#10000;
data_in <= 24'b011000110111101110010111;
#10000;
data_in <= 24'b011010011000000110011101;
#10000;
data_in <= 24'b011010000111111110011001;
#10000;
data_in <= 24'b010110110110111110001000;
#10000;
data_in <= 24'b011000110111101110010111;
#10000;
data_in <= 24'b011001011000000010011011;
#10000;
data_in <= 24'b011011011000010110100001;
#10000;
data_in <= 24'b011011111000011110100011;
#10000;
data_in <= 24'b011100101000101010100110;
#10000;
data_in <= 24'b011110101001000010101100;
#10000;
data_in <= 24'b011010111000000010011011;
#10000;
data_in <= 24'b010011010110000101111010;
#10000;
data_in <= 24'b010011100110010010000000;
#10000;
data_in <= 24'b010100110110101110000111;
#10000;
data_in <= 24'b011000000111011010010010;
#10000;
data_in <= 24'b011001010111101110010111;
#10000;
data_in <= 24'b011011001000001010011110;
#10000;
data_in <= 24'b011101101000110010101000;
#10000;
data_in <= 24'b011010111000000010011011;
#10000;
data_in <= 24'b010011110110001101111100;
#10000;
data_in <= 24'b001100100100100001100100;
#10000;
data_in <= 24'b001110100101000001101100;
#10000;
data_in <= 24'b010001000101101001110110;
#10000;
data_in <= 24'b010000010101011101110011;
#10000;
data_in <= 24'b001110100101000001101100;
#10000;
data_in <= 24'b001111010101001101101111;
#10000;
data_in <= 24'b001111010101001001101101;
#10000;
data_in <= 24'b001100010100010101011110;
#10000;
data_in <= 24'b001100000100010101100001;
#10000;
data_in <= 24'b001100010100011001100010;
#10000;
data_in <= 24'b001100110100100001100100;
#10000;
data_in <= 24'b001010010011111001011010;
#10000;
data_in <= 24'b000101110010110001001000;
#10000;
data_in <= 24'b000100010010011001000010;
#10000;
data_in <= 24'b000100110010011001000001;
#10000;
data_in <= 24'b000011000010000000111001;
#10000;
data_in <= 24'b001110000100110101101001;
#10000;
data_in <= 24'b001100000100010101100001;
#10000;
data_in <= 24'b001011100100001101011111;
#10000;
data_in <= 24'b001010110100000001011100;
#10000;
data_in <= 24'b000111110011010001010000;
#10000;
data_in <= 24'b000110000010110101001000;
#10000;
data_in <= 24'b000101000010011101000010;
#10000;
data_in <= 24'b000010100001111000110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101110100100001100010;
#10000;
data_in <= 24'b001100010011111101010101;
#10000;
data_in <= 24'b001001100011000001000010;
#10000;
data_in <= 24'b000110100010000100110000;
#10000;
data_in <= 24'b000101000001011000100001;
#10000;
data_in <= 24'b000011010000111100010111;
#10000;
data_in <= 24'b000011100000101100010100;
#10000;
data_in <= 24'b000011000000110000010010;
#10000;
data_in <= 24'b001111010100111001101000;
#10000;
data_in <= 24'b001011100011110001010010;
#10000;
data_in <= 24'b000111010010011100111001;
#10000;
data_in <= 24'b000100010001100000100111;
#10000;
data_in <= 24'b000010110000111100011010;
#10000;
data_in <= 24'b000001110000100000010010;
#10000;
data_in <= 24'b000001110000011000001111;
#10000;
data_in <= 24'b000010010000100100001111;
#10000;
data_in <= 24'b001111100100111101101001;
#10000;
data_in <= 24'b001010010011011101001101;
#10000;
data_in <= 24'b000101000001111100110011;
#10000;
data_in <= 24'b000011010001010100100110;
#10000;
data_in <= 24'b000010000000111000011011;
#10000;
data_in <= 24'b000000110000010100001111;
#10000;
data_in <= 24'b000000100000010000001100;
#10000;
data_in <= 24'b000001100000100000010000;
#10000;
data_in <= 24'b001101000100010101011111;
#10000;
data_in <= 24'b001000100011000001000110;
#10000;
data_in <= 24'b000100100001110100110001;
#10000;
data_in <= 24'b000011100001100000101001;
#10000;
data_in <= 24'b000010100001001000011111;
#10000;
data_in <= 24'b000000100000100000010011;
#10000;
data_in <= 24'b000001010000011100010001;
#10000;
data_in <= 24'b000010110001000000011001;
#10000;
data_in <= 24'b001000110011010001001110;
#10000;
data_in <= 24'b000101100010011100111100;
#10000;
data_in <= 24'b000010110001100100101100;
#10000;
data_in <= 24'b000010000001010000100110;
#10000;
data_in <= 24'b000001000000111100011101;
#10000;
data_in <= 24'b000000100000101100011000;
#10000;
data_in <= 24'b000011010001001100100000;
#10000;
data_in <= 24'b000110100010000000101101;
#10000;
data_in <= 24'b000100010010010100111110;
#10000;
data_in <= 24'b000010110001110100110100;
#10000;
data_in <= 24'b000001010001001100101001;
#10000;
data_in <= 24'b000000000000111000100001;
#10000;
data_in <= 24'b000000000000110100011101;
#10000;
data_in <= 24'b000001110001010000100010;
#10000;
data_in <= 24'b000110100010010100110011;
#10000;
data_in <= 24'b001010110011001101000100;
#10000;
data_in <= 24'b000001010001100100110010;
#10000;
data_in <= 24'b000010000001101000110001;
#10000;
data_in <= 24'b000001010001100000101101;
#10000;
data_in <= 24'b000001000001010100101000;
#10000;
data_in <= 24'b000011000001101100101110;
#10000;
data_in <= 24'b000110110010101100111100;
#10000;
data_in <= 24'b001010110011100101001011;
#10000;
data_in <= 24'b001100100100000001010010;
#10000;
data_in <= 24'b000000000001001100101100;
#10000;
data_in <= 24'b000001110001110000110010;
#10000;
data_in <= 24'b000011100010000000110111;
#10000;
data_in <= 24'b000100010010010000111001;
#10000;
data_in <= 24'b000111010011000001000101;
#10000;
data_in <= 24'b001100000100000101010100;
#10000;
data_in <= 24'b001101110100100001011011;
#10000;
data_in <= 24'b001101000100010101011010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000010110000111000010011;
#10000;
data_in <= 24'b000000110000011100001100;
#10000;
data_in <= 24'b000000110000100000001011;
#10000;
data_in <= 24'b000010100000111100010010;
#10000;
data_in <= 24'b000011100001001100010100;
#10000;
data_in <= 24'b000010010001000100010001;
#10000;
data_in <= 24'b000001110000111100001111;
#10000;
data_in <= 24'b000001100001001000010100;
#10000;
data_in <= 24'b000001010000100000010000;
#10000;
data_in <= 24'b000000100000100000001101;
#10000;
data_in <= 24'b000001100000101000001111;
#10000;
data_in <= 24'b000010000000111100010010;
#10000;
data_in <= 24'b000011000001000100010100;
#10000;
data_in <= 24'b000010100001000100010100;
#10000;
data_in <= 24'b000010100001001100010110;
#10000;
data_in <= 24'b000011000001100000011010;
#10000;
data_in <= 24'b000001000000100100010010;
#10000;
data_in <= 24'b000010000000111100011000;
#10000;
data_in <= 24'b000011010001001000011011;
#10000;
data_in <= 24'b000010110001001100011010;
#10000;
data_in <= 24'b000011010001001100011010;
#10000;
data_in <= 24'b000100000001100100011101;
#10000;
data_in <= 24'b000101100001111100100011;
#10000;
data_in <= 24'b000101010010000100100111;
#10000;
data_in <= 24'b000011110001010100100010;
#10000;
data_in <= 24'b000101010001110100101010;
#10000;
data_in <= 24'b000110010001111100101100;
#10000;
data_in <= 24'b000100110001110000100110;
#10000;
data_in <= 24'b000101010001111000101000;
#10000;
data_in <= 24'b000111100010011100110000;
#10000;
data_in <= 24'b001000110010110000110101;
#10000;
data_in <= 24'b001000010010101100110101;
#10000;
data_in <= 24'b001000000010011100111000;
#10000;
data_in <= 24'b001000100010101000111011;
#10000;
data_in <= 24'b001000100010100100111010;
#10000;
data_in <= 24'b000111100010011100110101;
#10000;
data_in <= 24'b001000110010110000111010;
#10000;
data_in <= 24'b001010100011010101000011;
#10000;
data_in <= 24'b001011000011011101000101;
#10000;
data_in <= 24'b001001010011001001000000;
#10000;
data_in <= 24'b001010100011001101000111;
#10000;
data_in <= 24'b001010010011000101001000;
#10000;
data_in <= 24'b001001110011000001000100;
#10000;
data_in <= 24'b001001110011000001000100;
#10000;
data_in <= 24'b001011000011011001001000;
#10000;
data_in <= 24'b001011110011101101001101;
#10000;
data_in <= 24'b001011110011101101001101;
#10000;
data_in <= 24'b001010010011011101001010;
#10000;
data_in <= 24'b001011010011011101001111;
#10000;
data_in <= 24'b001010110011010001001111;
#10000;
data_in <= 24'b001010110011010101001101;
#10000;
data_in <= 24'b001011110011100101010001;
#10000;
data_in <= 24'b001100010011101101010011;
#10000;
data_in <= 24'b001011100011101001010010;
#10000;
data_in <= 24'b001011110011101101010011;
#10000;
data_in <= 24'b001100000011111001010101;
#10000;
data_in <= 24'b001011000011100101010011;
#10000;
data_in <= 24'b001010100011011001010010;
#10000;
data_in <= 24'b001011010011100101010101;
#10000;
data_in <= 24'b001100110011111101011011;
#10000;
data_in <= 24'b001100110011111001011010;
#10000;
data_in <= 24'b001011000011100001010100;
#10000;
data_in <= 24'b001011110011101101010111;
#10000;
data_in <= 24'b001101010100001101011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000001010001000100010101;
#10000;
data_in <= 24'b000010010001100100100000;
#10000;
data_in <= 24'b000011110001111100101100;
#10000;
data_in <= 24'b000011110010000100110010;
#10000;
data_in <= 24'b000011110010000000111010;
#10000;
data_in <= 24'b000100000010010101000001;
#10000;
data_in <= 24'b000110000010110001001011;
#10000;
data_in <= 24'b000110010011001001010100;
#10000;
data_in <= 24'b000100010001110100100011;
#10000;
data_in <= 24'b000100110010001000101011;
#10000;
data_in <= 24'b000110000010011100110111;
#10000;
data_in <= 24'b000110010010101000111101;
#10000;
data_in <= 24'b000110000010110001000101;
#10000;
data_in <= 24'b000111010011001001001110;
#10000;
data_in <= 24'b001001100011101101011011;
#10000;
data_in <= 24'b001010100100001001100110;
#10000;
data_in <= 24'b000111000010100000110010;
#10000;
data_in <= 24'b000111000010110000111000;
#10000;
data_in <= 24'b001000000011000001000001;
#10000;
data_in <= 24'b001000010011001101001010;
#10000;
data_in <= 24'b001000110011100001010011;
#10000;
data_in <= 24'b001011000100000101100000;
#10000;
data_in <= 24'b001101110100110101110000;
#10000;
data_in <= 24'b001111100101100001111100;
#10000;
data_in <= 24'b001000100010111100111101;
#10000;
data_in <= 24'b001000010011000001000000;
#10000;
data_in <= 24'b001000100011001101001000;
#10000;
data_in <= 24'b001010000011100101010011;
#10000;
data_in <= 24'b001011010100000101100000;
#10000;
data_in <= 24'b001101110100111001101110;
#10000;
data_in <= 24'b010001010101110110000001;
#10000;
data_in <= 24'b010011110110101010001111;
#10000;
data_in <= 24'b001001100011010001000110;
#10000;
data_in <= 24'b001001000011001001001000;
#10000;
data_in <= 24'b001001010011011001010000;
#10000;
data_in <= 24'b001011010011111101011100;
#10000;
data_in <= 24'b001101110100110001101100;
#10000;
data_in <= 24'b010000110101100101111101;
#10000;
data_in <= 24'b010100110110101010010000;
#10000;
data_in <= 24'b011000000111101010100010;
#10000;
data_in <= 24'b001011010011101101010001;
#10000;
data_in <= 24'b001010100011100101010011;
#10000;
data_in <= 24'b001010110011110101011010;
#10000;
data_in <= 24'b001110000100101101101100;
#10000;
data_in <= 24'b010001000101101001111110;
#10000;
data_in <= 24'b010100000110011110001101;
#10000;
data_in <= 24'b011000010111101010100010;
#10000;
data_in <= 24'b011011101000101010110011;
#10000;
data_in <= 24'b001101000100001101011101;
#10000;
data_in <= 24'b001100000100000001011101;
#10000;
data_in <= 24'b001101000100100001100111;
#10000;
data_in <= 24'b010001000101100001111011;
#10000;
data_in <= 24'b010100010110100010001110;
#10000;
data_in <= 24'b010111010111011010011110;
#10000;
data_in <= 24'b011011101000011110110001;
#10000;
data_in <= 24'b011111001001011111000011;
#10000;
data_in <= 24'b001110000100100001100101;
#10000;
data_in <= 24'b001101000100011001100101;
#10000;
data_in <= 24'b001110010100110101110000;
#10000;
data_in <= 24'b010010100110000010000100;
#10000;
data_in <= 24'b010110100111000110010111;
#10000;
data_in <= 24'b011001010111111110100111;
#10000;
data_in <= 24'b011101001001000010111001;
#10000;
data_in <= 24'b100000101001111111001011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001010010100001101101011;
#10000;
data_in <= 24'b001100110101001101111100;
#10000;
data_in <= 24'b010001100110011010010001;
#10000;
data_in <= 24'b010011110111000110011100;
#10000;
data_in <= 24'b010101100111100110100101;
#10000;
data_in <= 24'b010111111000001010101110;
#10000;
data_in <= 24'b011001011000100110110111;
#10000;
data_in <= 24'b011010101000111010111100;
#10000;
data_in <= 24'b001101110101010001111011;
#10000;
data_in <= 24'b010000110110001110001100;
#10000;
data_in <= 24'b010100110111010110100000;
#10000;
data_in <= 24'b010111010111111110101010;
#10000;
data_in <= 24'b011000101000010110110001;
#10000;
data_in <= 24'b011001111000110010111000;
#10000;
data_in <= 24'b011011011001000110111111;
#10000;
data_in <= 24'b011011111001001111000001;
#10000;
data_in <= 24'b010011010110101010010001;
#10000;
data_in <= 24'b010110000111100010100001;
#10000;
data_in <= 24'b011001111000100110110100;
#10000;
data_in <= 24'b011011111001000110111100;
#10000;
data_in <= 24'b011100011001010011000000;
#10000;
data_in <= 24'b011100101001011011000100;
#10000;
data_in <= 24'b011101001001100011001000;
#10000;
data_in <= 24'b011100011001011111000111;
#10000;
data_in <= 24'b010111100111110010100101;
#10000;
data_in <= 24'b011001111000101010110010;
#10000;
data_in <= 24'b011101101001100011000011;
#10000;
data_in <= 24'b011110111001111011001010;
#10000;
data_in <= 24'b011110011001110111001011;
#10000;
data_in <= 24'b011101101001110111001010;
#10000;
data_in <= 24'b011101001001101011001010;
#10000;
data_in <= 24'b011100011001011111000111;
#10000;
data_in <= 24'b011011011000101110110100;
#10000;
data_in <= 24'b011101011001011111000010;
#10000;
data_in <= 24'b100000001010000111001110;
#10000;
data_in <= 24'b100000111010011011010010;
#10000;
data_in <= 24'b100000001010010011010010;
#10000;
data_in <= 24'b011110111010000111010001;
#10000;
data_in <= 24'b011101111001110011001110;
#10000;
data_in <= 24'b011100001001100011001001;
#10000;
data_in <= 24'b011110011001100111000100;
#10000;
data_in <= 24'b100000011010001111001110;
#10000;
data_in <= 24'b100010001010101111010111;
#10000;
data_in <= 24'b100001111010110011011000;
#10000;
data_in <= 24'b100001011010100111011001;
#10000;
data_in <= 24'b100000011010011111010111;
#10000;
data_in <= 24'b011110111010001111010100;
#10000;
data_in <= 24'b011101011001111011001111;
#10000;
data_in <= 24'b100001001010010011001111;
#10000;
data_in <= 24'b100010011010101111010110;
#10000;
data_in <= 24'b100011011011000011011100;
#10000;
data_in <= 24'b100010111011000011011100;
#10000;
data_in <= 24'b100010011010110111011101;
#10000;
data_in <= 24'b100001101010110011011100;
#10000;
data_in <= 24'b100000011010100111011010;
#10000;
data_in <= 24'b011111011010011011010111;
#10000;
data_in <= 24'b100010011010100111010100;
#10000;
data_in <= 24'b100011001010111011011001;
#10000;
data_in <= 24'b100011111011001011011101;
#10000;
data_in <= 24'b100011001011000111011101;
#10000;
data_in <= 24'b100010111010111111011101;
#10000;
data_in <= 24'b100001111010111111011111;
#10000;
data_in <= 24'b100001011010110111011110;
#10000;
data_in <= 24'b100000011010101011011011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000101000011010110110;
#10000;
data_in <= 24'b011001101000101010111010;
#10000;
data_in <= 24'b011001101000101010111000;
#10000;
data_in <= 24'b011000011000010110110011;
#10000;
data_in <= 24'b011000001000000110101110;
#10000;
data_in <= 24'b010111000111110110101010;
#10000;
data_in <= 24'b010101100111100010100011;
#10000;
data_in <= 24'b010100000111000010011011;
#10000;
data_in <= 24'b011010101000111010111110;
#10000;
data_in <= 24'b011011011001000111000001;
#10000;
data_in <= 24'b011011011001000111000001;
#10000;
data_in <= 24'b011010001000110010111010;
#10000;
data_in <= 24'b011001101000100010110110;
#10000;
data_in <= 24'b011001101000011110110100;
#10000;
data_in <= 24'b011000101000001110110000;
#10000;
data_in <= 24'b010111000111111010101001;
#10000;
data_in <= 24'b011010111001000011000010;
#10000;
data_in <= 24'b011011001001001011000010;
#10000;
data_in <= 24'b011010101001000011000000;
#10000;
data_in <= 24'b011010001000110010111010;
#10000;
data_in <= 24'b011001101000101010111000;
#10000;
data_in <= 24'b011010001000101110110111;
#10000;
data_in <= 24'b011001111000101010110110;
#10000;
data_in <= 24'b011001011000011010110011;
#10000;
data_in <= 24'b011011101001001111000101;
#10000;
data_in <= 24'b011011011001001011000100;
#10000;
data_in <= 24'b011010011000111011000000;
#10000;
data_in <= 24'b011001011000101110111011;
#10000;
data_in <= 24'b011001011000100110111001;
#10000;
data_in <= 24'b011001011000100110110111;
#10000;
data_in <= 24'b011001011000100110110111;
#10000;
data_in <= 24'b011001111000101010110110;
#10000;
data_in <= 24'b011101001001101111001111;
#10000;
data_in <= 24'b011100011001100111001010;
#10000;
data_in <= 24'b011011001001010011000101;
#10000;
data_in <= 24'b011010001001000011000000;
#10000;
data_in <= 24'b011001111000110110111101;
#10000;
data_in <= 24'b011001011000110010111001;
#10000;
data_in <= 24'b011001011000110010111001;
#10000;
data_in <= 24'b011010001000110010111010;
#10000;
data_in <= 24'b011110001010000011010100;
#10000;
data_in <= 24'b011100111001101111001111;
#10000;
data_in <= 24'b011011111001100011001001;
#10000;
data_in <= 24'b011011011001010111000110;
#10000;
data_in <= 24'b011010011001000111000010;
#10000;
data_in <= 24'b011001101000110010111100;
#10000;
data_in <= 24'b011001011000101110111011;
#10000;
data_in <= 24'b011001101000110010111100;
#10000;
data_in <= 24'b011110011010000111010101;
#10000;
data_in <= 24'b011100101001110111010000;
#10000;
data_in <= 24'b011011111001101011001101;
#10000;
data_in <= 24'b011100001001100111001010;
#10000;
data_in <= 24'b011010111001010011000101;
#10000;
data_in <= 24'b011001011000110110111110;
#10000;
data_in <= 24'b011000101000101010111011;
#10000;
data_in <= 24'b011000111000101110111100;
#10000;
data_in <= 24'b011110101010010111011000;
#10000;
data_in <= 24'b011101011010000011010011;
#10000;
data_in <= 24'b011100111001111011010001;
#10000;
data_in <= 24'b011100111001111011010001;
#10000;
data_in <= 24'b011100011001101011001011;
#10000;
data_in <= 24'b011010011001001011000011;
#10000;
data_in <= 24'b011001101000111010111111;
#10000;
data_in <= 24'b011001101000111111000000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010101000111000110011101;
#10000;
data_in <= 24'b010011110110101010010110;
#10000;
data_in <= 24'b010001100101111110001001;
#10000;
data_in <= 24'b001111000101010101111111;
#10000;
data_in <= 24'b001110100101001101111011;
#10000;
data_in <= 24'b001110010101001101111000;
#10000;
data_in <= 24'b001101100100110101110011;
#10000;
data_in <= 24'b001011100100011101101001;
#10000;
data_in <= 24'b011000100111111110101011;
#10000;
data_in <= 24'b010111110111101010100110;
#10000;
data_in <= 24'b010101110111001010011110;
#10000;
data_in <= 24'b010100010110101010010100;
#10000;
data_in <= 24'b010011110110100010010010;
#10000;
data_in <= 24'b010011100110011110001111;
#10000;
data_in <= 24'b010001110110000110000110;
#10000;
data_in <= 24'b010000010101100101111101;
#10000;
data_in <= 24'b011010111000101010110111;
#10000;
data_in <= 24'b011010111000100010110100;
#10000;
data_in <= 24'b011001111000010010110000;
#10000;
data_in <= 24'b011000101000000010101001;
#10000;
data_in <= 24'b011000110111111110101000;
#10000;
data_in <= 24'b011000110111110110100101;
#10000;
data_in <= 24'b010110110111010110011101;
#10000;
data_in <= 24'b010100110110110110010010;
#10000;
data_in <= 24'b011010111000110010111001;
#10000;
data_in <= 24'b011010101000101110111000;
#10000;
data_in <= 24'b011001111000100010110101;
#10000;
data_in <= 24'b011001101000011010110001;
#10000;
data_in <= 24'b011001111000010010110000;
#10000;
data_in <= 24'b011001101000010010101101;
#10000;
data_in <= 24'b011000100111111010100111;
#10000;
data_in <= 24'b010110110111100010011111;
#10000;
data_in <= 24'b011001101000101010111000;
#10000;
data_in <= 24'b011010001000101010111000;
#10000;
data_in <= 24'b011001001000011010110100;
#10000;
data_in <= 24'b011000001000001110101111;
#10000;
data_in <= 24'b011000001000000110101110;
#10000;
data_in <= 24'b011000101000010010101111;
#10000;
data_in <= 24'b011000011000000110101100;
#10000;
data_in <= 24'b010111000111110010100101;
#10000;
data_in <= 24'b011001001000101010111010;
#10000;
data_in <= 24'b011001001000101010111010;
#10000;
data_in <= 24'b011000001000011010110110;
#10000;
data_in <= 24'b010110111000001010101111;
#10000;
data_in <= 24'b010111001000000010101110;
#10000;
data_in <= 24'b010111111000010010110000;
#10000;
data_in <= 24'b011000001000001110101111;
#10000;
data_in <= 24'b010111101000000010101011;
#10000;
data_in <= 24'b011000101000101010111011;
#10000;
data_in <= 24'b011000101000101010111011;
#10000;
data_in <= 24'b010111111000011110111000;
#10000;
data_in <= 24'b010110101000001010110010;
#10000;
data_in <= 24'b010110111000000110110001;
#10000;
data_in <= 24'b010111011000010010110001;
#10000;
data_in <= 24'b010111111000001110110001;
#10000;
data_in <= 24'b010111001000000110101101;
#10000;
data_in <= 24'b010111111000100010111001;
#10000;
data_in <= 24'b011000001000100110111010;
#10000;
data_in <= 24'b010111101000011110111000;
#10000;
data_in <= 24'b010110101000001110110100;
#10000;
data_in <= 24'b010110011000000110110010;
#10000;
data_in <= 24'b010110101000001010110010;
#10000;
data_in <= 24'b010110111000000110110001;
#10000;
data_in <= 24'b010110000111111110101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101110100101101101110;
#10000;
data_in <= 24'b001111110101010001110100;
#10000;
data_in <= 24'b010000000101001001110001;
#10000;
data_in <= 24'b001101100100100001100111;
#10000;
data_in <= 24'b001101000100010001100001;
#10000;
data_in <= 24'b001101010100010101100010;
#10000;
data_in <= 24'b001011010011101101010111;
#10000;
data_in <= 24'b000111000010101001000110;
#10000;
data_in <= 24'b001101110100110101110000;
#10000;
data_in <= 24'b001110100100111101101111;
#10000;
data_in <= 24'b001101100100100101101010;
#10000;
data_in <= 24'b001011010100000101100000;
#10000;
data_in <= 24'b001011000011111001011101;
#10000;
data_in <= 24'b001011100100000001011101;
#10000;
data_in <= 24'b001010110011101101011000;
#10000;
data_in <= 24'b001000100011001101001110;
#10000;
data_in <= 24'b010000100101101001111110;
#10000;
data_in <= 24'b001111000101001001110101;
#10000;
data_in <= 24'b001100100100100101101001;
#10000;
data_in <= 24'b001010110100000001011111;
#10000;
data_in <= 24'b001001110011101101011010;
#10000;
data_in <= 24'b001001000011100001010111;
#10000;
data_in <= 24'b001000110011010101010100;
#10000;
data_in <= 24'b001000010011001101010000;
#10000;
data_in <= 24'b010101100111000010010101;
#10000;
data_in <= 24'b010010000110001010000110;
#10000;
data_in <= 24'b001111010101011001111000;
#10000;
data_in <= 24'b001101010100111001101110;
#10000;
data_in <= 24'b001011000100001101100011;
#10000;
data_in <= 24'b000111110011011001010110;
#10000;
data_in <= 24'b000110100010111101001111;
#10000;
data_in <= 24'b000110100010111001001101;
#10000;
data_in <= 24'b010111110111110010100011;
#10000;
data_in <= 24'b010100110111000010010101;
#10000;
data_in <= 24'b010010110110011010001011;
#10000;
data_in <= 24'b010001110110001110000110;
#10000;
data_in <= 24'b001111000101011001111010;
#10000;
data_in <= 24'b001010010100010001100110;
#10000;
data_in <= 24'b000111010011011001011000;
#10000;
data_in <= 24'b000111010011010001010100;
#10000;
data_in <= 24'b010110110111101110100100;
#10000;
data_in <= 24'b010101010111011010011101;
#10000;
data_in <= 24'b010100110111001010011001;
#10000;
data_in <= 24'b010100110111001110010111;
#10000;
data_in <= 24'b010011000110100110001110;
#10000;
data_in <= 24'b001111000101100101111110;
#10000;
data_in <= 24'b001011110100101001101111;
#10000;
data_in <= 24'b001011010100011001101000;
#10000;
data_in <= 24'b010110100111110110101001;
#10000;
data_in <= 24'b010110000111101110100110;
#10000;
data_in <= 24'b010101110111100110100100;
#10000;
data_in <= 24'b010101010111100010100000;
#10000;
data_in <= 24'b010100010111000110011010;
#10000;
data_in <= 24'b010001110110100010001111;
#10000;
data_in <= 24'b001111010101110010000011;
#10000;
data_in <= 24'b001110010101010001111001;
#10000;
data_in <= 24'b010111011000000110101111;
#10000;
data_in <= 24'b010111001000000110101101;
#10000;
data_in <= 24'b010110100111110110101001;
#10000;
data_in <= 24'b010101000111011110100010;
#10000;
data_in <= 24'b010011110111001010011101;
#10000;
data_in <= 24'b010010010110110010010100;
#10000;
data_in <= 24'b001111110110000110001100;
#10000;
data_in <= 24'b001111000101100110000000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000011100001110000111000;
#10000;
data_in <= 24'b000010010001100000110010;
#10000;
data_in <= 24'b000010000001011000101101;
#10000;
data_in <= 24'b000011000001101100101110;
#10000;
data_in <= 24'b000101110010001100110101;
#10000;
data_in <= 24'b000111100010101100111001;
#10000;
data_in <= 24'b001000110010110100110111;
#10000;
data_in <= 24'b001000010010110000110100;
#10000;
data_in <= 24'b000110110010100101000101;
#10000;
data_in <= 24'b000101000010001100111101;
#10000;
data_in <= 24'b000011010001101100110010;
#10000;
data_in <= 24'b000010100001100000101011;
#10000;
data_in <= 24'b000011000001100000101010;
#10000;
data_in <= 24'b000011100001100100100111;
#10000;
data_in <= 24'b000011110001100100100011;
#10000;
data_in <= 24'b000011010001100000100000;
#10000;
data_in <= 24'b001000000011000101001100;
#10000;
data_in <= 24'b000110110010101001000100;
#10000;
data_in <= 24'b000101000010001000111001;
#10000;
data_in <= 24'b000011010001101100101110;
#10000;
data_in <= 24'b000010100001011100100111;
#10000;
data_in <= 24'b000010100001011000100010;
#10000;
data_in <= 24'b000010100001010000011110;
#10000;
data_in <= 24'b000010110001010000011101;
#10000;
data_in <= 24'b000111010010110101001010;
#10000;
data_in <= 24'b000111000010101101000101;
#10000;
data_in <= 24'b000110010010011100111110;
#10000;
data_in <= 24'b000101000010001000110101;
#10000;
data_in <= 24'b000100000001110100101101;
#10000;
data_in <= 24'b000011100001101000100110;
#10000;
data_in <= 24'b000011100001011100100001;
#10000;
data_in <= 24'b000011010001011100011110;
#10000;
data_in <= 24'b000111000010110001001001;
#10000;
data_in <= 24'b000111010010110001000110;
#10000;
data_in <= 24'b000111000010101001000001;
#10000;
data_in <= 24'b000110000010011000111001;
#10000;
data_in <= 24'b000100100001111100101111;
#10000;
data_in <= 24'b000011000001100000100100;
#10000;
data_in <= 24'b000010000001000100011010;
#10000;
data_in <= 24'b000001000000111000010101;
#10000;
data_in <= 24'b000111110011000101010000;
#10000;
data_in <= 24'b001000000010111101001001;
#10000;
data_in <= 24'b000110110010101101000010;
#10000;
data_in <= 24'b000110000010011100111010;
#10000;
data_in <= 24'b000101010010001000110010;
#10000;
data_in <= 24'b000100000001110000101000;
#10000;
data_in <= 24'b000010110001011000011110;
#10000;
data_in <= 24'b000001110001000100011000;
#10000;
data_in <= 24'b001010010011111001011101;
#10000;
data_in <= 24'b001001010011011001010001;
#10000;
data_in <= 24'b000111000010101101000101;
#10000;
data_in <= 24'b000101100010010000111010;
#10000;
data_in <= 24'b000101100010001000110100;
#10000;
data_in <= 24'b000101100010000100101111;
#10000;
data_in <= 24'b000101010001111100101001;
#10000;
data_in <= 24'b000100110001110100100100;
#10000;
data_in <= 24'b001101110100111001101110;
#10000;
data_in <= 24'b001011010011111101011100;
#10000;
data_in <= 24'b000110110010110001000111;
#10000;
data_in <= 24'b000011110001111100110110;
#10000;
data_in <= 24'b000011100001110000101111;
#10000;
data_in <= 24'b000100000001110100101011;
#10000;
data_in <= 24'b000101000001111000101000;
#10000;
data_in <= 24'b000101000001111000100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000101100010000000100111;
#10000;
data_in <= 24'b000110110010010100101100;
#10000;
data_in <= 24'b000111000010010100101110;
#10000;
data_in <= 24'b000101000001110100100110;
#10000;
data_in <= 24'b000010010001001100011101;
#10000;
data_in <= 24'b000010010001001100011101;
#10000;
data_in <= 24'b000101000001110100101011;
#10000;
data_in <= 24'b000111110010100000110101;
#10000;
data_in <= 24'b000101010001111100100110;
#10000;
data_in <= 24'b000110010010001100101010;
#10000;
data_in <= 24'b000111000010010100101110;
#10000;
data_in <= 24'b000101110010000000101001;
#10000;
data_in <= 24'b000100000001100100100011;
#10000;
data_in <= 24'b000011110001100100100011;
#10000;
data_in <= 24'b000101110010000000101101;
#10000;
data_in <= 24'b001000010010100100110110;
#10000;
data_in <= 24'b000101000001110000100011;
#10000;
data_in <= 24'b000110000010000100100101;
#10000;
data_in <= 24'b000110110010001100101010;
#10000;
data_in <= 24'b000101110010000100101000;
#10000;
data_in <= 24'b000101000001110100100110;
#10000;
data_in <= 24'b000100110001110000100110;
#10000;
data_in <= 24'b000101100001111000101011;
#10000;
data_in <= 24'b000110100010001100101101;
#10000;
data_in <= 24'b000011110001100000011100;
#10000;
data_in <= 24'b000100010001101000011110;
#10000;
data_in <= 24'b000100110001110000100000;
#10000;
data_in <= 24'b000101000001110000100011;
#10000;
data_in <= 24'b000100110001101100100010;
#10000;
data_in <= 24'b000100000001100100100010;
#10000;
data_in <= 24'b000100010001011100100010;
#10000;
data_in <= 24'b000100010001011100100010;
#10000;
data_in <= 24'b000010000001000100010101;
#10000;
data_in <= 24'b000010110001001000010101;
#10000;
data_in <= 24'b000011000001001100010110;
#10000;
data_in <= 24'b000011110001010100011010;
#10000;
data_in <= 24'b000100010001011100011110;
#10000;
data_in <= 24'b000100000001011100100000;
#10000;
data_in <= 24'b000100000001010100011110;
#10000;
data_in <= 24'b000011010001010000011101;
#10000;
data_in <= 24'b000001110000110100010010;
#10000;
data_in <= 24'b000001110000111000010001;
#10000;
data_in <= 24'b000010000000111100010010;
#10000;
data_in <= 24'b000010110001001000010101;
#10000;
data_in <= 24'b000011110001010100011010;
#10000;
data_in <= 24'b000100100001100000011111;
#10000;
data_in <= 24'b000100110001100100100000;
#10000;
data_in <= 24'b000101000001101000100001;
#10000;
data_in <= 24'b000010110001000100010110;
#10000;
data_in <= 24'b000010100001000100010100;
#10000;
data_in <= 24'b000010100000111100010010;
#10000;
data_in <= 24'b000010100000111100010010;
#10000;
data_in <= 24'b000011010001001000010101;
#10000;
data_in <= 24'b000100010001010100011010;
#10000;
data_in <= 24'b000101010001100100011110;
#10000;
data_in <= 24'b000101100001110000100011;
#10000;
data_in <= 24'b000100000001100100011101;
#10000;
data_in <= 24'b000011110001011000011001;
#10000;
data_in <= 24'b000011010001001000010101;
#10000;
data_in <= 24'b000010010000111000010001;
#10000;
data_in <= 24'b000010010000111000010001;
#10000;
data_in <= 24'b000011000001000100010100;
#10000;
data_in <= 24'b000100100001011000011011;
#10000;
data_in <= 24'b000101100001101000011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001000110010101000110011;
#10000;
data_in <= 24'b000110000010000000100111;
#10000;
data_in <= 24'b000111010010010100101100;
#10000;
data_in <= 24'b001100100011101001000001;
#10000;
data_in <= 24'b001101110011110101000010;
#10000;
data_in <= 24'b001001110010110100110010;
#10000;
data_in <= 24'b001000110010100000101011;
#10000;
data_in <= 24'b001010100010111100110010;
#10000;
data_in <= 24'b001001010010110000110101;
#10000;
data_in <= 24'b000111010010010100101100;
#10000;
data_in <= 24'b001000010010100100110000;
#10000;
data_in <= 24'b001100010011100101000000;
#10000;
data_in <= 24'b001101010011101101000000;
#10000;
data_in <= 24'b001001110010110100110010;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b001001010010101000101101;
#10000;
data_in <= 24'b001000110010101000110011;
#10000;
data_in <= 24'b001000010010100100110000;
#10000;
data_in <= 24'b001001010010110100110100;
#10000;
data_in <= 24'b001011110011011100111110;
#10000;
data_in <= 24'b001100100011100000111101;
#10000;
data_in <= 24'b001010010010111100110100;
#10000;
data_in <= 24'b001000110010100000101011;
#10000;
data_in <= 24'b001000000010010100101000;
#10000;
data_in <= 24'b000110100010000100101010;
#10000;
data_in <= 24'b000111000010010000101011;
#10000;
data_in <= 24'b001000100010101000110001;
#10000;
data_in <= 24'b001010010011000100111000;
#10000;
data_in <= 24'b001011110011010100111010;
#10000;
data_in <= 24'b001011000011001000110111;
#10000;
data_in <= 24'b001001110010110000101111;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b000011000001010000011011;
#10000;
data_in <= 24'b000100010001100100100000;
#10000;
data_in <= 24'b000110000010000000100111;
#10000;
data_in <= 24'b001000000010100000101111;
#10000;
data_in <= 24'b001010010010111100110100;
#10000;
data_in <= 24'b001010110011000100110110;
#10000;
data_in <= 24'b001010010010111000110001;
#10000;
data_in <= 24'b001001000010100100101100;
#10000;
data_in <= 24'b000001100000111000010101;
#10000;
data_in <= 24'b000010000001000000010111;
#10000;
data_in <= 24'b000011110001011100011110;
#10000;
data_in <= 24'b000110010010000100101000;
#10000;
data_in <= 24'b001001000010101000101111;
#10000;
data_in <= 24'b001001100010110000110001;
#10000;
data_in <= 24'b001001110010110000101111;
#10000;
data_in <= 24'b001001010010101000101101;
#10000;
data_in <= 24'b000011110001011100011110;
#10000;
data_in <= 24'b000011000001010000011011;
#10000;
data_in <= 24'b000100000001100000011111;
#10000;
data_in <= 24'b000110110010001100101010;
#10000;
data_in <= 24'b001001010010101100110000;
#10000;
data_in <= 24'b001001000010101000101111;
#10000;
data_in <= 24'b001001010010101000101101;
#10000;
data_in <= 24'b001001110010110000101111;
#10000;
data_in <= 24'b000111010010001100101010;
#10000;
data_in <= 24'b000101000001110000100011;
#10000;
data_in <= 24'b000101100001111000100101;
#10000;
data_in <= 24'b001000010010100100110000;
#10000;
data_in <= 24'b001010000010111000110011;
#10000;
data_in <= 24'b001001000010101000101111;
#10000;
data_in <= 24'b001001010010101000101101;
#10000;
data_in <= 24'b001010010010111000110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001000010010010100100110;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001010010010101100101011;
#10000;
data_in <= 24'b001010010010101100101011;
#10000;
data_in <= 24'b001011010010111100101111;
#10000;
data_in <= 24'b001100100011010000110100;
#10000;
data_in <= 24'b001100010011001000110000;
#10000;
data_in <= 24'b001010110010110000101010;
#10000;
data_in <= 24'b001000010010010100100110;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001010100010110000101100;
#10000;
data_in <= 24'b001011100011000000110000;
#10000;
data_in <= 24'b001011100010111100101101;
#10000;
data_in <= 24'b001010010010101000101000;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010010010101100101011;
#10000;
data_in <= 24'b001011010010111100101111;
#10000;
data_in <= 24'b001011100010111100101101;
#10000;
data_in <= 24'b001011000010110100101011;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001010000010101000101010;
#10000;
data_in <= 24'b001010110010110100101101;
#10000;
data_in <= 24'b001011110011000000101110;
#10000;
data_in <= 24'b001011110011000000101110;
#10000;
data_in <= 24'b001000010010010100100110;
#10000;
data_in <= 24'b001000010010010100100110;
#10000;
data_in <= 24'b001000110010010100100101;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010100010110000101100;
#10000;
data_in <= 24'b001011110011000000101110;
#10000;
data_in <= 24'b001100100011001100110001;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001010000010101000101010;
#10000;
data_in <= 24'b001010110010110100101101;
#10000;
data_in <= 24'b001011000010111000101110;
#10000;
data_in <= 24'b001011010010111100101111;
#10000;
data_in <= 24'b001100110011010000110010;
#10000;
data_in <= 24'b001110000011100100110111;
#10000;
data_in <= 24'b001010010010110100101110;
#10000;
data_in <= 24'b001010000010110000101101;
#10000;
data_in <= 24'b001011000010111000101110;
#10000;
data_in <= 24'b001100000011001000110010;
#10000;
data_in <= 24'b001011110011000100110001;
#10000;
data_in <= 24'b001011100011000000110000;
#10000;
data_in <= 24'b001100110011010000110010;
#10000;
data_in <= 24'b001110000011100100110111;
#10000;
data_in <= 24'b001001110010101100101100;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001010010010101100101011;
#10000;
data_in <= 24'b001011000010111000101110;
#10000;
data_in <= 24'b001010110010110100101101;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010110010110000101010;
#10000;
data_in <= 24'b001100010011001000110000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000110111100010010111;
#10000;
data_in <= 24'b010100010110011010000101;
#10000;
data_in <= 24'b001110100100111101101011;
#10000;
data_in <= 24'b001011010100001001011110;
#10000;
data_in <= 24'b001011110100010001011111;
#10000;
data_in <= 24'b001100110100100001100011;
#10000;
data_in <= 24'b001011010100000001011011;
#10000;
data_in <= 24'b001000000011010001001101;
#10000;
data_in <= 24'b010110110111000010001111;
#10000;
data_in <= 24'b010100100110011110000110;
#10000;
data_in <= 24'b010010100101111101111011;
#10000;
data_in <= 24'b010010100101111101111011;
#10000;
data_in <= 24'b010101000110100110000100;
#10000;
data_in <= 24'b010110110111000010001011;
#10000;
data_in <= 24'b010101000110100010000001;
#10000;
data_in <= 24'b010001110101101101110100;
#10000;
data_in <= 24'b010100010110100110000111;
#10000;
data_in <= 24'b010100000110100010000110;
#10000;
data_in <= 24'b010101000110101010000110;
#10000;
data_in <= 24'b010111000111001010001110;
#10000;
data_in <= 24'b011010000111110110011000;
#10000;
data_in <= 24'b011010100111111110011010;
#10000;
data_in <= 24'b010111100111001010001011;
#10000;
data_in <= 24'b010011110110001101111100;
#10000;
data_in <= 24'b010011010110010110000011;
#10000;
data_in <= 24'b010011010110010110000011;
#10000;
data_in <= 24'b010100000110100010000100;
#10000;
data_in <= 24'b010110010110111110001011;
#10000;
data_in <= 24'b010111100111010110001111;
#10000;
data_in <= 24'b010110010110111010001001;
#10000;
data_in <= 24'b010010100101111001110111;
#10000;
data_in <= 24'b001110110100111101101000;
#10000;
data_in <= 24'b010100010110101110001001;
#10000;
data_in <= 24'b010011100110100010000110;
#10000;
data_in <= 24'b010011000110011110000010;
#10000;
data_in <= 24'b010011110110011110000011;
#10000;
data_in <= 24'b010100010110100010000010;
#10000;
data_in <= 24'b010010100101111101111010;
#10000;
data_in <= 24'b010000000101010001101101;
#10000;
data_in <= 24'b001101110100101101100100;
#10000;
data_in <= 24'b010111100111101010011000;
#10000;
data_in <= 24'b010101010111000110001111;
#10000;
data_in <= 24'b010011000110100110000100;
#10000;
data_in <= 24'b010001110110001001111101;
#10000;
data_in <= 24'b010000110101110001110110;
#10000;
data_in <= 24'b001111010101010001101110;
#10000;
data_in <= 24'b001101110100110101100110;
#10000;
data_in <= 24'b001101110100101101100100;
#10000;
data_in <= 24'b011000111000000110011110;
#10000;
data_in <= 24'b010101100111010010010001;
#10000;
data_in <= 24'b010010000110010110000000;
#10000;
data_in <= 24'b001111010101100001110011;
#10000;
data_in <= 24'b001100110100110001100110;
#10000;
data_in <= 24'b001010100100000101011011;
#10000;
data_in <= 24'b001001110011110101010110;
#10000;
data_in <= 24'b001010010011111101011000;
#10000;
data_in <= 24'b010111000111101010010101;
#10000;
data_in <= 24'b010100000110110110001000;
#10000;
data_in <= 24'b010000100101110101111000;
#10000;
data_in <= 24'b001101010100111001101000;
#10000;
data_in <= 24'b001010010100000001011010;
#10000;
data_in <= 24'b000111100011010101001111;
#10000;
data_in <= 24'b000111000011000101001100;
#10000;
data_in <= 24'b001000000011010101010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000101110010101101000100;
#10000;
data_in <= 24'b000101000010100100111111;
#10000;
data_in <= 24'b000110010010111001000100;
#10000;
data_in <= 24'b001001010011101001010000;
#10000;
data_in <= 24'b001010100011111101010101;
#10000;
data_in <= 24'b001010000011101101010000;
#10000;
data_in <= 24'b001010000011101101010000;
#10000;
data_in <= 24'b001011010011111101010110;
#10000;
data_in <= 24'b010000010101010101101110;
#10000;
data_in <= 24'b001100000100010001011101;
#10000;
data_in <= 24'b001001010011100101010010;
#10000;
data_in <= 24'b001011000100000001011001;
#10000;
data_in <= 24'b001101100100101001100011;
#10000;
data_in <= 24'b001101010100100101100010;
#10000;
data_in <= 24'b001011110100001101011100;
#10000;
data_in <= 24'b001010110011111001011001;
#10000;
data_in <= 24'b010010110101111101111000;
#10000;
data_in <= 24'b001110100100111001100111;
#10000;
data_in <= 24'b001011100100010001011101;
#10000;
data_in <= 24'b001101000100100101100100;
#10000;
data_in <= 24'b001111100101001101101110;
#10000;
data_in <= 24'b001111010101001001101101;
#10000;
data_in <= 24'b001101100100101101100110;
#10000;
data_in <= 24'b001100000100010101100001;
#10000;
data_in <= 24'b001101100100101001100011;
#10000;
data_in <= 24'b001110010100110101100110;
#10000;
data_in <= 24'b001111100101001101101110;
#10000;
data_in <= 24'b010001010101101001110110;
#10000;
data_in <= 24'b010001000101100101110101;
#10000;
data_in <= 24'b001110110101000001101111;
#10000;
data_in <= 24'b001101110100110001101011;
#10000;
data_in <= 24'b001110000100110101101100;
#10000;
data_in <= 24'b001100110100011101100000;
#10000;
data_in <= 24'b010000010101010101101110;
#10000;
data_in <= 24'b010011110110010001111111;
#10000;
data_in <= 24'b010101000110100110000101;
#10000;
data_in <= 24'b010010100101111101111110;
#10000;
data_in <= 24'b001111010101001001110010;
#10000;
data_in <= 24'b001110000100110101101101;
#10000;
data_in <= 24'b001110110101000001110000;
#10000;
data_in <= 24'b001110010100110101100110;
#10000;
data_in <= 24'b010000110101011101110000;
#10000;
data_in <= 24'b010011110110010010000000;
#10000;
data_in <= 24'b010101000110100010000111;
#10000;
data_in <= 24'b010011100110001110000011;
#10000;
data_in <= 24'b010001010101101001111010;
#10000;
data_in <= 24'b001111010101001101110110;
#10000;
data_in <= 24'b001111100101001001110101;
#10000;
data_in <= 24'b001101010100100101100010;
#10000;
data_in <= 24'b010000010101010101101110;
#10000;
data_in <= 24'b010100000110001001111111;
#10000;
data_in <= 24'b010101000110100010000111;
#10000;
data_in <= 24'b010011110110010010000100;
#10000;
data_in <= 24'b010010000101110001111111;
#10000;
data_in <= 24'b010000000101011001111010;
#10000;
data_in <= 24'b001111110101001101110110;
#10000;
data_in <= 24'b001100000100010101100000;
#10000;
data_in <= 24'b010001010101101001110101;
#10000;
data_in <= 24'b010110010110111010001010;
#10000;
data_in <= 24'b010111010111000110010000;
#10000;
data_in <= 24'b010100000110010010000111;
#10000;
data_in <= 24'b010000110101011101111010;
#10000;
data_in <= 24'b001111010101000001110101;
#10000;
data_in <= 24'b001111100101000101110100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001100010011111101011011;
#10000;
data_in <= 24'b001100110100000101011110;
#10000;
data_in <= 24'b001101010100001101100000;
#10000;
data_in <= 24'b001110000100011001100011;
#10000;
data_in <= 24'b001111000100011101100101;
#10000;
data_in <= 24'b001110110100100101100110;
#10000;
data_in <= 24'b001110110100100101100110;
#10000;
data_in <= 24'b001110010100100001101000;
#10000;
data_in <= 24'b001101000100011001100011;
#10000;
data_in <= 24'b001101110100011001100110;
#10000;
data_in <= 24'b001110110100100001101000;
#10000;
data_in <= 24'b001111010100101001101010;
#10000;
data_in <= 24'b001111110100110001101100;
#10000;
data_in <= 24'b010000010100111001101110;
#10000;
data_in <= 24'b010000000100111101101111;
#10000;
data_in <= 24'b001111100101000001101111;
#10000;
data_in <= 24'b001110100100110001101011;
#10000;
data_in <= 24'b001110100100101101101100;
#10000;
data_in <= 24'b001111010100110001101101;
#10000;
data_in <= 24'b001111110100111001101111;
#10000;
data_in <= 24'b010000010101000001110001;
#10000;
data_in <= 24'b010001000101001101110100;
#10000;
data_in <= 24'b010001100101010101110110;
#10000;
data_in <= 24'b010001010101011001110111;
#10000;
data_in <= 24'b001110010100110001101101;
#10000;
data_in <= 24'b001111000100110101101110;
#10000;
data_in <= 24'b001111100100110101101110;
#10000;
data_in <= 24'b010000000100111101110000;
#10000;
data_in <= 24'b010000100101000101110010;
#10000;
data_in <= 24'b010001010101010001110101;
#10000;
data_in <= 24'b010010000101011101111000;
#10000;
data_in <= 24'b010001110101100001111001;
#10000;
data_in <= 24'b001110100100110101101110;
#10000;
data_in <= 24'b001111010100111101101110;
#10000;
data_in <= 24'b001111110100111001101110;
#10000;
data_in <= 24'b010000010101000001110000;
#10000;
data_in <= 24'b010001000101001101110100;
#10000;
data_in <= 24'b010001110101011001110111;
#10000;
data_in <= 24'b010010100101100101111010;
#10000;
data_in <= 24'b010010010101101001111011;
#10000;
data_in <= 24'b001111010101000101110000;
#10000;
data_in <= 24'b010000000101001001110001;
#10000;
data_in <= 24'b010000110101001001110010;
#10000;
data_in <= 24'b010001010101010001110100;
#10000;
data_in <= 24'b010010000101011101111000;
#10000;
data_in <= 24'b010010110101101001111011;
#10000;
data_in <= 24'b010011010101110001111101;
#10000;
data_in <= 24'b010011110101111001111111;
#10000;
data_in <= 24'b001111110101001101110010;
#10000;
data_in <= 24'b010000100101010001110001;
#10000;
data_in <= 24'b010001110101011101110100;
#10000;
data_in <= 24'b010010100101101001110111;
#10000;
data_in <= 24'b010011010101110001111100;
#10000;
data_in <= 24'b010011110101111001111110;
#10000;
data_in <= 24'b010100010110000010000000;
#10000;
data_in <= 24'b010100100110000110000001;
#10000;
data_in <= 24'b010000010101001101110010;
#10000;
data_in <= 24'b010001010101010101110010;
#10000;
data_in <= 24'b010010000101100001110101;
#10000;
data_in <= 24'b010011000101110001111001;
#10000;
data_in <= 24'b010011110101111001111110;
#10000;
data_in <= 24'b010100010110000010000000;
#10000;
data_in <= 24'b010100100110000110000001;
#10000;
data_in <= 24'b010100100110000110000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001110000100101001101001;
#10000;
data_in <= 24'b001110000100101101101100;
#10000;
data_in <= 24'b010000110101011101111010;
#10000;
data_in <= 24'b010101000110110010010000;
#10000;
data_in <= 24'b011001111000000110100110;
#10000;
data_in <= 24'b011101111001000110111001;
#10000;
data_in <= 24'b100001001010000011001001;
#10000;
data_in <= 24'b100011011010101111010100;
#10000;
data_in <= 24'b001111010100111001101111;
#10000;
data_in <= 24'b001111110101001101110110;
#10000;
data_in <= 24'b010011100110000110000110;
#10000;
data_in <= 24'b011000010111100110011101;
#10000;
data_in <= 24'b011101001000111010110011;
#10000;
data_in <= 24'b100000011001101111000011;
#10000;
data_in <= 24'b100011001010100111010000;
#10000;
data_in <= 24'b100100101011000111011000;
#10000;
data_in <= 24'b010000110101001101110111;
#10000;
data_in <= 24'b010010010101110110000000;
#10000;
data_in <= 24'b010111000110111110010100;
#10000;
data_in <= 24'b011100001000100010101100;
#10000;
data_in <= 24'b100000101001110011000000;
#10000;
data_in <= 24'b100011101010100111001110;
#10000;
data_in <= 24'b100101011011001011010111;
#10000;
data_in <= 24'b100110011011100111011101;
#10000;
data_in <= 24'b010010000101100001111100;
#10000;
data_in <= 24'b010100010110010110001000;
#10000;
data_in <= 24'b011001100111101010011101;
#10000;
data_in <= 24'b011110101001001110110101;
#10000;
data_in <= 24'b100010111010010111001001;
#10000;
data_in <= 24'b100101101011001011010101;
#10000;
data_in <= 24'b100111101011101011011101;
#10000;
data_in <= 24'b101000001011111011100001;
#10000;
data_in <= 24'b010011110110000010000001;
#10000;
data_in <= 24'b010110100110111110001111;
#10000;
data_in <= 24'b011011111000010010100100;
#10000;
data_in <= 24'b100000011001101010111010;
#10000;
data_in <= 24'b100100011010110011001110;
#10000;
data_in <= 24'b100111011011100111011011;
#10000;
data_in <= 24'b101001101100001011100100;
#10000;
data_in <= 24'b101010011100010111100111;
#10000;
data_in <= 24'b010101100110011110001000;
#10000;
data_in <= 24'b011001000111011110011000;
#10000;
data_in <= 24'b011110011000111010101110;
#10000;
data_in <= 24'b100010111010001011000010;
#10000;
data_in <= 24'b100110101011001111010011;
#10000;
data_in <= 24'b101001101100001011100000;
#10000;
data_in <= 24'b101011101100101111101010;
#10000;
data_in <= 24'b101100011100111011101101;
#10000;
data_in <= 24'b010110010110101110001010;
#10000;
data_in <= 24'b011010100111111010011101;
#10000;
data_in <= 24'b100000011001011010110101;
#10000;
data_in <= 24'b100100111010101111001001;
#10000;
data_in <= 24'b101000011011101111011001;
#10000;
data_in <= 24'b101011011100101011100101;
#10000;
data_in <= 24'b101100111101000111101110;
#10000;
data_in <= 24'b101101001101001011101111;
#10000;
data_in <= 24'b010110010110101110001010;
#10000;
data_in <= 24'b011011001000000010011111;
#10000;
data_in <= 24'b100001101001101010111001;
#10000;
data_in <= 24'b100110101010111111001110;
#10000;
data_in <= 24'b101001111011111111011101;
#10000;
data_in <= 24'b101100101100110111101000;
#10000;
data_in <= 24'b101101011101000111101111;
#10000;
data_in <= 24'b101101011101000111101111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100101011011010111011110;
#10000;
data_in <= 24'b100100111011011011011110;
#10000;
data_in <= 24'b100100101011010111100000;
#10000;
data_in <= 24'b100011111011010011100000;
#10000;
data_in <= 24'b100011101011001011100000;
#10000;
data_in <= 24'b100001111010111111011111;
#10000;
data_in <= 24'b100001011010110111011110;
#10000;
data_in <= 24'b100000111010110011011101;
#10000;
data_in <= 24'b100110111011101011100001;
#10000;
data_in <= 24'b100110011011101011100001;
#10000;
data_in <= 24'b100101111011101011100010;
#10000;
data_in <= 24'b100101011011100011100011;
#10000;
data_in <= 24'b100100011011011011100010;
#10000;
data_in <= 24'b100011001011001111100000;
#10000;
data_in <= 24'b100010001011000011100000;
#10000;
data_in <= 24'b100001101010111111100000;
#10000;
data_in <= 24'b101000011100000111100101;
#10000;
data_in <= 24'b100111111100000111100101;
#10000;
data_in <= 24'b100111101011111111100110;
#10000;
data_in <= 24'b100110101011110111100101;
#10000;
data_in <= 24'b100101011011101111100101;
#10000;
data_in <= 24'b100100001011011111100011;
#10000;
data_in <= 24'b100011001011010111100010;
#10000;
data_in <= 24'b100010011011001111100010;
#10000;
data_in <= 24'b101010011100011111101010;
#10000;
data_in <= 24'b101001101100011011101001;
#10000;
data_in <= 24'b101001001100010011101000;
#10000;
data_in <= 24'b100111111100000011100111;
#10000;
data_in <= 24'b100110101011111011100110;
#10000;
data_in <= 24'b100101011011101111100101;
#10000;
data_in <= 24'b100100011011100011100100;
#10000;
data_in <= 24'b100011011011011011100011;
#10000;
data_in <= 24'b101011101100101011101100;
#10000;
data_in <= 24'b101010101100100111101010;
#10000;
data_in <= 24'b101010001100011011101001;
#10000;
data_in <= 24'b101000111100001111100111;
#10000;
data_in <= 24'b100111001100000011100110;
#10000;
data_in <= 24'b100110001011110011100100;
#10000;
data_in <= 24'b100101001011101011100100;
#10000;
data_in <= 24'b100100011011100011100100;
#10000;
data_in <= 24'b101011111100110011101011;
#10000;
data_in <= 24'b101011101100101111101010;
#10000;
data_in <= 24'b101010111100011111101001;
#10000;
data_in <= 24'b101001001100010011100111;
#10000;
data_in <= 24'b100111111100000111100101;
#10000;
data_in <= 24'b100110101011111011100100;
#10000;
data_in <= 24'b100110001011110011100100;
#10000;
data_in <= 24'b100101011011101111100101;
#10000;
data_in <= 24'b101100011100110111101011;
#10000;
data_in <= 24'b101011111100110011101011;
#10000;
data_in <= 24'b101011001100100111101000;
#10000;
data_in <= 24'b101001111100011011100111;
#10000;
data_in <= 24'b101000101100001011100110;
#10000;
data_in <= 24'b100111001100000011100110;
#10000;
data_in <= 24'b100110101011111011100110;
#10000;
data_in <= 24'b100110001011111011101000;
#10000;
data_in <= 24'b101100101100111011101100;
#10000;
data_in <= 24'b101100001100110011101010;
#10000;
data_in <= 24'b101011001100100111101000;
#10000;
data_in <= 24'b101001111100011011100101;
#10000;
data_in <= 24'b101000111100010011100101;
#10000;
data_in <= 24'b100111111100001011100100;
#10000;
data_in <= 24'b100111011100000111100101;
#10000;
data_in <= 24'b100111001100000011100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011111101010100111011100;
#10000;
data_in <= 24'b011110011010010011010111;
#10000;
data_in <= 24'b011101001001111111010010;
#10000;
data_in <= 24'b011100011001110011001111;
#10000;
data_in <= 24'b011100001001101111001100;
#10000;
data_in <= 24'b011011101001100111001010;
#10000;
data_in <= 24'b011010111001010011000101;
#10000;
data_in <= 24'b011001111001000011000001;
#10000;
data_in <= 24'b100001001010110111011110;
#10000;
data_in <= 24'b011111011010100011011011;
#10000;
data_in <= 24'b011101111010001011010101;
#10000;
data_in <= 24'b011101001001111111010010;
#10000;
data_in <= 24'b011100111001111011001111;
#10000;
data_in <= 24'b011100011001110011001101;
#10000;
data_in <= 24'b011011101001011111001000;
#10000;
data_in <= 24'b011010101001001111000100;
#10000;
data_in <= 24'b100010001011000111100010;
#10000;
data_in <= 24'b100001001010110111011110;
#10000;
data_in <= 24'b011111001010011111011000;
#10000;
data_in <= 24'b011110011010010011010101;
#10000;
data_in <= 24'b011110011010001011010011;
#10000;
data_in <= 24'b011101101001111111010000;
#10000;
data_in <= 24'b011100101001110011001011;
#10000;
data_in <= 24'b011011101001011111001000;
#10000;
data_in <= 24'b100010111011001111100011;
#10000;
data_in <= 24'b100001111011000011100001;
#10000;
data_in <= 24'b100000101010101111011100;
#10000;
data_in <= 24'b011111001010011111011000;
#10000;
data_in <= 24'b011111001010010111010110;
#10000;
data_in <= 24'b011110011010001111010010;
#10000;
data_in <= 24'b011101011001111111001110;
#10000;
data_in <= 24'b011100111001101111001011;
#10000;
data_in <= 24'b100011001011010111100010;
#10000;
data_in <= 24'b100010011011001111100010;
#10000;
data_in <= 24'b100001011010111111011110;
#10000;
data_in <= 24'b100000101010110011011011;
#10000;
data_in <= 24'b100000001010100011011000;
#10000;
data_in <= 24'b011111101010011111010100;
#10000;
data_in <= 24'b011110111010010011010001;
#10000;
data_in <= 24'b011110011010000111010001;
#10000;
data_in <= 24'b100100001011011111100011;
#10000;
data_in <= 24'b100011011011011011100011;
#10000;
data_in <= 24'b100010111011001111100011;
#10000;
data_in <= 24'b100010001011001011100001;
#10000;
data_in <= 24'b100001101010111111011100;
#10000;
data_in <= 24'b100001001010110111011010;
#10000;
data_in <= 24'b100000111010110011011001;
#10000;
data_in <= 24'b100001011010110011011001;
#10000;
data_in <= 24'b100101001011101111100111;
#10000;
data_in <= 24'b100100101011110011100111;
#10000;
data_in <= 24'b100100011011101011100111;
#10000;
data_in <= 24'b100100001011100111100110;
#10000;
data_in <= 24'b100011101011011111100100;
#10000;
data_in <= 24'b100011011011011011100011;
#10000;
data_in <= 24'b100011111011011011100010;
#10000;
data_in <= 24'b100100001011011111100100;
#10000;
data_in <= 24'b100110111011111111100111;
#10000;
data_in <= 24'b100110101100000111101000;
#10000;
data_in <= 24'b100110001100000011101010;
#10000;
data_in <= 24'b100101111011111111101001;
#10000;
data_in <= 24'b100101101011111011101000;
#10000;
data_in <= 24'b100101101011111011101000;
#10000;
data_in <= 24'b100101111011111111101001;
#10000;
data_in <= 24'b100110101100000011101010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011001111000111111000011;
#10000;
data_in <= 24'b011001001000111111000010;
#10000;
data_in <= 24'b011000111000101110111111;
#10000;
data_in <= 24'b011000001000100110111010;
#10000;
data_in <= 24'b010111101000011110111000;
#10000;
data_in <= 24'b010111001000011010110101;
#10000;
data_in <= 24'b010111001000010010110100;
#10000;
data_in <= 24'b010111001000010110110010;
#10000;
data_in <= 24'b011001111000111111000011;
#10000;
data_in <= 24'b011001111000111111000011;
#10000;
data_in <= 24'b011001101000111011000010;
#10000;
data_in <= 24'b011001011000110111000001;
#10000;
data_in <= 24'b011001001000110110111110;
#10000;
data_in <= 24'b011000101000101110111100;
#10000;
data_in <= 24'b011000101000101010111010;
#10000;
data_in <= 24'b011000011000100110111001;
#10000;
data_in <= 24'b011100011001100111001101;
#10000;
data_in <= 24'b011100001001011111001011;
#10000;
data_in <= 24'b011011011001010111000110;
#10000;
data_in <= 24'b011010011001000111000010;
#10000;
data_in <= 24'b011001111000111111000000;
#10000;
data_in <= 24'b011001011000110110111110;
#10000;
data_in <= 24'b011001111000110010111110;
#10000;
data_in <= 24'b011001111000110110111101;
#10000;
data_in <= 24'b011110001010000011010001;
#10000;
data_in <= 24'b011101011001110011010000;
#10000;
data_in <= 24'b011100101001011111001001;
#10000;
data_in <= 24'b011011001001010011000101;
#10000;
data_in <= 24'b011010111001000011000010;
#10000;
data_in <= 24'b011011001001000111000011;
#10000;
data_in <= 24'b011011101001001111000101;
#10000;
data_in <= 24'b011011111001010011000110;
#10000;
data_in <= 24'b011110001001110111001111;
#10000;
data_in <= 24'b011110001001110111001111;
#10000;
data_in <= 24'b011110101001110111001111;
#10000;
data_in <= 24'b011101111001110011001110;
#10000;
data_in <= 24'b011101111001101111001011;
#10000;
data_in <= 24'b011101101001101011001010;
#10000;
data_in <= 24'b011101001001100011001000;
#10000;
data_in <= 24'b011100111001011111000111;
#10000;
data_in <= 24'b100001001010100011011000;
#10000;
data_in <= 24'b100001011010100011011010;
#10000;
data_in <= 24'b100001101010100111011011;
#10000;
data_in <= 24'b100000111010011011011000;
#10000;
data_in <= 24'b011111101001111111010000;
#10000;
data_in <= 24'b011100111001010011000101;
#10000;
data_in <= 24'b011010011000101010111011;
#10000;
data_in <= 24'b011000101000001110110100;
#10000;
data_in <= 24'b100101001011100011101000;
#10000;
data_in <= 24'b100100101011001111100100;
#10000;
data_in <= 24'b100010101010101111011100;
#10000;
data_in <= 24'b011111111010000011010001;
#10000;
data_in <= 24'b011100101001001011000011;
#10000;
data_in <= 24'b011001011000010110110110;
#10000;
data_in <= 24'b010110010111100110101010;
#10000;
data_in <= 24'b010100110111001110100100;
#10000;
data_in <= 24'b100110101011110011101010;
#10000;
data_in <= 24'b100100001011001011100000;
#10000;
data_in <= 24'b100000011010001011010000;
#10000;
data_in <= 24'b011100001001000110111111;
#10000;
data_in <= 24'b011000101000001110110001;
#10000;
data_in <= 24'b010110100111101110101001;
#10000;
data_in <= 24'b010101110111011110101000;
#10000;
data_in <= 24'b010101100111011110100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010111111000011010110011;
#10000;
data_in <= 24'b010111101000010110110010;
#10000;
data_in <= 24'b010111101000001010110000;
#10000;
data_in <= 24'b010110100111111110101011;
#10000;
data_in <= 24'b010101000111100110100101;
#10000;
data_in <= 24'b010011110111001010011101;
#10000;
data_in <= 24'b010010010110110010011000;
#10000;
data_in <= 24'b010010010110100110010010;
#10000;
data_in <= 24'b011000111000100110111001;
#10000;
data_in <= 24'b011000001000011110110100;
#10000;
data_in <= 24'b010111101000001010110000;
#10000;
data_in <= 24'b010110010111110110101011;
#10000;
data_in <= 24'b010100110111100010100100;
#10000;
data_in <= 24'b010011010111001010011110;
#10000;
data_in <= 24'b010001110110110010011000;
#10000;
data_in <= 24'b010001110110100110010100;
#10000;
data_in <= 24'b011010001000111010111110;
#10000;
data_in <= 24'b011001011000101110111011;
#10000;
data_in <= 24'b011001001000100010110110;
#10000;
data_in <= 24'b011000011000010110110011;
#10000;
data_in <= 24'b010111101000001010110000;
#10000;
data_in <= 24'b010101110111101110101001;
#10000;
data_in <= 24'b010011110111001110100001;
#10000;
data_in <= 24'b010011000110110110011010;
#10000;
data_in <= 24'b011011011001000111000001;
#10000;
data_in <= 24'b011010111000111110111111;
#10000;
data_in <= 24'b011010001000110010111010;
#10000;
data_in <= 24'b011001111000101110111001;
#10000;
data_in <= 24'b011000111000011110110101;
#10000;
data_in <= 24'b010110110111111110101101;
#10000;
data_in <= 24'b010100000111010010100010;
#10000;
data_in <= 24'b010010110110110010011001;
#10000;
data_in <= 24'b011100101001001111000100;
#10000;
data_in <= 24'b011011111001000011000001;
#10000;
data_in <= 24'b011010111000110110111011;
#10000;
data_in <= 24'b011010001000101010111000;
#10000;
data_in <= 24'b011001011000011110110101;
#10000;
data_in <= 24'b011000011000001110110001;
#10000;
data_in <= 24'b010110110111110110101011;
#10000;
data_in <= 24'b010110000111100110100111;
#10000;
data_in <= 24'b010110000111100110101010;
#10000;
data_in <= 24'b010101100111011110101000;
#10000;
data_in <= 24'b010100110111010110100011;
#10000;
data_in <= 24'b010100010111001110100001;
#10000;
data_in <= 24'b010100110111010110100011;
#10000;
data_in <= 24'b010101110111100110100111;
#10000;
data_in <= 24'b010111010111111110101101;
#10000;
data_in <= 24'b011000101000001110110001;
#10000;
data_in <= 24'b010001010110011010010100;
#10000;
data_in <= 24'b010010000110100110010111;
#10000;
data_in <= 24'b010010110110110010011010;
#10000;
data_in <= 24'b010010100110101110011001;
#10000;
data_in <= 24'b010010010110101010011000;
#10000;
data_in <= 24'b010010100110101110011001;
#10000;
data_in <= 24'b010011010110111010011100;
#10000;
data_in <= 24'b010100010111001010100000;
#10000;
data_in <= 24'b011010001000100110110111;
#10000;
data_in <= 24'b011011111001000010111110;
#10000;
data_in <= 24'b011101011001011011000100;
#10000;
data_in <= 24'b011100101001001111000000;
#10000;
data_in <= 24'b011001101000011110110100;
#10000;
data_in <= 24'b010110010111101010100111;
#10000;
data_in <= 24'b010100010111000010011101;
#10000;
data_in <= 24'b010011100110110010011011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010001000101110010000000;
#10000;
data_in <= 24'b001100110100011101100110;
#10000;
data_in <= 24'b000111110011000101001110;
#10000;
data_in <= 24'b000101110010100001000010;
#10000;
data_in <= 24'b000100110010000100110111;
#10000;
data_in <= 24'b000010100001100100101001;
#10000;
data_in <= 24'b000010100001011000100010;
#10000;
data_in <= 24'b000011110001100000100001;
#10000;
data_in <= 24'b010010010110001110001000;
#10000;
data_in <= 24'b010000100101011001111001;
#10000;
data_in <= 24'b001011010100000001100001;
#10000;
data_in <= 24'b000110100010110101001000;
#10000;
data_in <= 24'b000100000010000000110111;
#10000;
data_in <= 24'b000011000001110000101101;
#10000;
data_in <= 24'b000011010001100000100110;
#10000;
data_in <= 24'b000010110001010100011111;
#10000;
data_in <= 24'b010011110110100110010001;
#10000;
data_in <= 24'b010011100110011010001010;
#10000;
data_in <= 24'b001111000101001001110101;
#10000;
data_in <= 24'b001000100011011001010101;
#10000;
data_in <= 24'b000100110010010000111110;
#10000;
data_in <= 24'b000100000010000100110100;
#10000;
data_in <= 24'b000100010001111000101110;
#10000;
data_in <= 24'b000010110001011100100011;
#10000;
data_in <= 24'b010100000110101110010111;
#10000;
data_in <= 24'b010100010110101010010010;
#10000;
data_in <= 24'b010001100101110110000011;
#10000;
data_in <= 24'b001100000100011101100111;
#10000;
data_in <= 24'b000111010011001001001101;
#10000;
data_in <= 24'b000101010010100000111101;
#10000;
data_in <= 24'b000100100010001000110011;
#10000;
data_in <= 24'b000011110001110100101001;
#10000;
data_in <= 24'b010100110111000010011101;
#10000;
data_in <= 24'b010011100110101010010011;
#10000;
data_in <= 24'b010010000110001010001010;
#10000;
data_in <= 24'b010000000101100001111100;
#10000;
data_in <= 24'b001011110100010001100011;
#10000;
data_in <= 24'b000110110010111101001000;
#10000;
data_in <= 24'b000100010010001000110101;
#10000;
data_in <= 24'b000100010010000100101110;
#10000;
data_in <= 24'b010101110111010110100100;
#10000;
data_in <= 24'b010011110110110010011001;
#10000;
data_in <= 24'b010010110110011110010000;
#10000;
data_in <= 24'b010010100110010110001010;
#10000;
data_in <= 24'b001111110101011001110110;
#10000;
data_in <= 24'b001001100011101101010110;
#10000;
data_in <= 24'b000101010010100000111101;
#10000;
data_in <= 24'b000100110010001100110011;
#10000;
data_in <= 24'b010110010111011110100110;
#10000;
data_in <= 24'b010100100111000010011111;
#10000;
data_in <= 24'b010011100110101110010111;
#10000;
data_in <= 24'b010011000110100110010000;
#10000;
data_in <= 24'b010010000110000110000011;
#10000;
data_in <= 24'b001110010100111101101011;
#10000;
data_in <= 24'b001001000011100101001111;
#10000;
data_in <= 24'b000101110010100100111010;
#10000;
data_in <= 24'b010101010111011010100100;
#10000;
data_in <= 24'b010100110111010010100010;
#10000;
data_in <= 24'b010011100110110110011010;
#10000;
data_in <= 24'b010010110110011110010000;
#10000;
data_in <= 24'b010010100110011010001001;
#10000;
data_in <= 24'b010001100101111101111111;
#10000;
data_in <= 24'b001100100100011101100010;
#10000;
data_in <= 24'b000111010011000001000101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000100110001101100100010;
#10000;
data_in <= 24'b000100110001100100011110;
#10000;
data_in <= 24'b000101000001100100011100;
#10000;
data_in <= 24'b000100100001011100011010;
#10000;
data_in <= 24'b000011100001000100010101;
#10000;
data_in <= 24'b000010000000101100001111;
#10000;
data_in <= 24'b000001110000101000001111;
#10000;
data_in <= 24'b000010100000111000010011;
#10000;
data_in <= 24'b000100010001101100100010;
#10000;
data_in <= 24'b000011100001011100011011;
#10000;
data_in <= 24'b000011110001010100011010;
#10000;
data_in <= 24'b000101000001100100011100;
#10000;
data_in <= 24'b000101110001101000011110;
#10000;
data_in <= 24'b000101000001011100011011;
#10000;
data_in <= 24'b000100010001010000011001;
#10000;
data_in <= 24'b000100000001010000011001;
#10000;
data_in <= 24'b000011110001100000100001;
#10000;
data_in <= 24'b000010010001001000010110;
#10000;
data_in <= 24'b000010000000111000010011;
#10000;
data_in <= 24'b000100000001011000011011;
#10000;
data_in <= 24'b000111000010000000100101;
#10000;
data_in <= 24'b000111110010001100101000;
#10000;
data_in <= 24'b000111010010000100100110;
#10000;
data_in <= 24'b000110100001111000100011;
#10000;
data_in <= 24'b000011010001011100100001;
#10000;
data_in <= 24'b000001000000111000010101;
#10000;
data_in <= 24'b000000000000100000001111;
#10000;
data_in <= 24'b000010000000111000010011;
#10000;
data_in <= 24'b000100110001100100011110;
#10000;
data_in <= 24'b000111000010000000100101;
#10000;
data_in <= 24'b001000000010010000101001;
#10000;
data_in <= 24'b001000000010011000101011;
#10000;
data_in <= 24'b000100000001110000101000;
#10000;
data_in <= 24'b000010000001001100011011;
#10000;
data_in <= 24'b000000000000101000010001;
#10000;
data_in <= 24'b000000000000100000001111;
#10000;
data_in <= 24'b000001000000101000010001;
#10000;
data_in <= 24'b000010100001000000010111;
#10000;
data_in <= 24'b000100110001100100100000;
#10000;
data_in <= 24'b000110110010000100101000;
#10000;
data_in <= 24'b000101100010010000110000;
#10000;
data_in <= 24'b000100000001110000100110;
#10000;
data_in <= 24'b000010000001001100011011;
#10000;
data_in <= 24'b000000010000101100010010;
#10000;
data_in <= 24'b000000000000010000001011;
#10000;
data_in <= 24'b000000000000001100001010;
#10000;
data_in <= 24'b000001000000101000010001;
#10000;
data_in <= 24'b000011010001001100011010;
#10000;
data_in <= 24'b000101010010010100110010;
#10000;
data_in <= 24'b000101010010000100101011;
#10000;
data_in <= 24'b000100010001110000100100;
#10000;
data_in <= 24'b000011000001010100011110;
#10000;
data_in <= 24'b000001010000110000010101;
#10000;
data_in <= 24'b000000000000010100001110;
#10000;
data_in <= 24'b000000000000010100001110;
#10000;
data_in <= 24'b000000100000100100010010;
#10000;
data_in <= 24'b000100010010000100110010;
#10000;
data_in <= 24'b000100000010000000101101;
#10000;
data_in <= 24'b000101000010000000101010;
#10000;
data_in <= 24'b000101010010000000101000;
#10000;
data_in <= 24'b000100000001100100100010;
#10000;
data_in <= 24'b000010000000111100011000;
#10000;
data_in <= 24'b000000010000100100010000;
#10000;
data_in <= 24'b000000000000100000001111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000100010001011100011110;
#10000;
data_in <= 24'b000011000001010000011011;
#10000;
data_in <= 24'b000011100001011000011101;
#10000;
data_in <= 24'b000110010010000100101000;
#10000;
data_in <= 24'b001000110010100100101110;
#10000;
data_in <= 24'b001001010010101100110000;
#10000;
data_in <= 24'b001001110010110000101111;
#10000;
data_in <= 24'b001010000010110100110000;
#10000;
data_in <= 24'b000100000001011000011101;
#10000;
data_in <= 24'b000010110001001100011010;
#10000;
data_in <= 24'b000011010001010100011100;
#10000;
data_in <= 24'b000101100001111000100101;
#10000;
data_in <= 24'b000111110010010100101010;
#10000;
data_in <= 24'b001000000010011000101011;
#10000;
data_in <= 24'b001000000010010100101000;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b000011010001001100011010;
#10000;
data_in <= 24'b000010010001000100011000;
#10000;
data_in <= 24'b000011000001010000011011;
#10000;
data_in <= 24'b000101000001110000100011;
#10000;
data_in <= 24'b000111010010001100101000;
#10000;
data_in <= 24'b000111110010010100101010;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b000100110001101100100010;
#10000;
data_in <= 24'b000100100001101000100001;
#10000;
data_in <= 24'b000100100001101000100001;
#10000;
data_in <= 24'b000101010001110100100100;
#10000;
data_in <= 24'b000110110010000100100110;
#10000;
data_in <= 24'b000111100010010000101001;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b000111100010011000101101;
#10000;
data_in <= 24'b000111000010010000101011;
#10000;
data_in <= 24'b000110000010000000100111;
#10000;
data_in <= 24'b000101100001111000100101;
#10000;
data_in <= 24'b000110000001111000100011;
#10000;
data_in <= 24'b000110100010000000100101;
#10000;
data_in <= 24'b000111010010001000100101;
#10000;
data_in <= 24'b000111010010001000100101;
#10000;
data_in <= 24'b000100110001101100100010;
#10000;
data_in <= 24'b000101010001110100100100;
#10000;
data_in <= 24'b000101000001110000100011;
#10000;
data_in <= 24'b000100100001101000100001;
#10000;
data_in <= 24'b000101100001110000100001;
#10000;
data_in <= 24'b000111000010001000100111;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b000000110000101100010010;
#10000;
data_in <= 24'b000010010001000100011000;
#10000;
data_in <= 24'b000011110001011100011110;
#10000;
data_in <= 24'b000100010001100100100000;
#10000;
data_in <= 24'b000110000001111000100011;
#10000;
data_in <= 24'b000111110010010100101010;
#10000;
data_in <= 24'b001001000010100100101100;
#10000;
data_in <= 24'b001000110010100000101011;
#10000;
data_in <= 24'b000000100000101000010001;
#10000;
data_in <= 24'b000010100001001000011001;
#10000;
data_in <= 24'b000100100001101000100001;
#10000;
data_in <= 24'b000101000001110000100011;
#10000;
data_in <= 24'b000101110010000000100100;
#10000;
data_in <= 24'b000110110010010000101000;
#10000;
data_in <= 24'b000111000010001100100110;
#10000;
data_in <= 24'b000110000001111100100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001001100010101000101011;
#10000;
data_in <= 24'b001001100010101000101011;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010010010101000101000;
#10000;
data_in <= 24'b001010010010101000101000;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001001010010100100101010;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010010010101000101000;
#10000;
data_in <= 24'b001010100010101100101001;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010100010101100101001;
#10000;
data_in <= 24'b001010110010110000101010;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010100010101100101001;
#10000;
data_in <= 24'b001010110010110000101010;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001001110010100100101001;
#10000;
data_in <= 24'b001010100010101100101001;
#10000;
data_in <= 24'b001010110010110000101010;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001100010100000101000;
#10000;
data_in <= 24'b001010010010101000101000;
#10000;
data_in <= 24'b001010100010101100101001;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001010000010100100100111;
#10000;
data_in <= 24'b001010000010100100100111;
#10000;
data_in <= 24'b001000110010100000101001;
#10000;
data_in <= 24'b001000110010100000101001;
#10000;
data_in <= 24'b001000110010100000100111;
#10000;
data_in <= 24'b001000110010100000100111;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001010010100000100110;
#10000;
data_in <= 24'b001001110010100000100110;
#10000;
data_in <= 24'b001010000010100100100111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010001100110000101111011;
#10000;
data_in <= 24'b010010110110010001111110;
#10000;
data_in <= 24'b010010000101111101111001;
#10000;
data_in <= 24'b001101010100101001100101;
#10000;
data_in <= 24'b001000010011010001001111;
#10000;
data_in <= 24'b000110000010101101000110;
#10000;
data_in <= 24'b000110110011000001001011;
#10000;
data_in <= 24'b001000100011100001010100;
#10000;
data_in <= 24'b010110110111010110001101;
#10000;
data_in <= 24'b010100110110101110000011;
#10000;
data_in <= 24'b010001010101100101110010;
#10000;
data_in <= 24'b001101000100010101011111;
#10000;
data_in <= 24'b001001000011001001001110;
#10000;
data_in <= 24'b000110110010110001000111;
#10000;
data_in <= 24'b001000010011001101010000;
#10000;
data_in <= 24'b001010100100000001011100;
#10000;
data_in <= 24'b011000010111100110010001;
#10000;
data_in <= 24'b010010010110000101111001;
#10000;
data_in <= 24'b001100110100011101100000;
#10000;
data_in <= 24'b001001110011100001010010;
#10000;
data_in <= 24'b001000000010111001001010;
#10000;
data_in <= 24'b000111000010110101001000;
#10000;
data_in <= 24'b001001110011100101010110;
#10000;
data_in <= 24'b001101110100110101101001;
#10000;
data_in <= 24'b010100010110011110000000;
#10000;
data_in <= 24'b001101100100110001100101;
#10000;
data_in <= 24'b001001000011010101001111;
#10000;
data_in <= 24'b001000010011001001001100;
#10000;
data_in <= 24'b001000100011000001001100;
#10000;
data_in <= 24'b001000010011001001001101;
#10000;
data_in <= 24'b001100010100001101100000;
#10000;
data_in <= 24'b010001110101110001111011;
#10000;
data_in <= 24'b010001000101100001110001;
#10000;
data_in <= 24'b001100000100000101011011;
#10000;
data_in <= 24'b001000110011010001001110;
#10000;
data_in <= 24'b001010000011011101010001;
#10000;
data_in <= 24'b001010000011011001010010;
#10000;
data_in <= 24'b001001100011011001010011;
#10000;
data_in <= 24'b001110000100101001101001;
#10000;
data_in <= 24'b010100100110011110000110;
#10000;
data_in <= 24'b010000110101010001101110;
#10000;
data_in <= 24'b001100010100001001011100;
#10000;
data_in <= 24'b001010000011011101010001;
#10000;
data_in <= 24'b001010000011011001010010;
#10000;
data_in <= 24'b001001100011010001010001;
#10000;
data_in <= 24'b001001010011010001010100;
#10000;
data_in <= 24'b001110010100101101101010;
#10000;
data_in <= 24'b010100000110011110000111;
#10000;
data_in <= 24'b010011000101110001110011;
#10000;
data_in <= 24'b001110010100100001100010;
#10000;
data_in <= 24'b001010100011011101010001;
#10000;
data_in <= 24'b001001000011000001001100;
#10000;
data_in <= 24'b001000100011000001001101;
#10000;
data_in <= 24'b001010000011011101010111;
#10000;
data_in <= 24'b001111100101000101110010;
#10000;
data_in <= 24'b010101110110110110010000;
#10000;
data_in <= 24'b010101010110010101111100;
#10000;
data_in <= 24'b001111110100111101100110;
#10000;
data_in <= 24'b001010100011011001010010;
#10000;
data_in <= 24'b001000010010110101001001;
#10000;
data_in <= 24'b001000100010111101001111;
#10000;
data_in <= 24'b001100100100000101100010;
#10000;
data_in <= 24'b010011100110000110000100;
#10000;
data_in <= 24'b011001010111111010100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001111010101001101101111;
#10000;
data_in <= 24'b010110010111000110001111;
#10000;
data_in <= 24'b011000100111101110011011;
#10000;
data_in <= 24'b010101110110110110010000;
#10000;
data_in <= 24'b010011010110000110000100;
#10000;
data_in <= 24'b010010000101101001111111;
#10000;
data_in <= 24'b010001100101010101111100;
#10000;
data_in <= 24'b010010100101011101111101;
#10000;
data_in <= 24'b010001110101111101111101;
#10000;
data_in <= 24'b010110110111011110010110;
#10000;
data_in <= 24'b011000000111101110011101;
#10000;
data_in <= 24'b010011110110101010001100;
#10000;
data_in <= 24'b010001110101110110000001;
#10000;
data_in <= 24'b010001100101100001111101;
#10000;
data_in <= 24'b010010010101010101111101;
#10000;
data_in <= 24'b010011110101101010000000;
#10000;
data_in <= 24'b010101000110111010001100;
#10000;
data_in <= 24'b011000100111111010011101;
#10000;
data_in <= 24'b010111100111100110011011;
#10000;
data_in <= 24'b010010100110010110000111;
#10000;
data_in <= 24'b010000110101100101111101;
#10000;
data_in <= 24'b010000110101011001111100;
#10000;
data_in <= 24'b010010000101011101111110;
#10000;
data_in <= 24'b010100100101110110000011;
#10000;
data_in <= 24'b010111100111011110010111;
#10000;
data_in <= 24'b011001001000000110100000;
#10000;
data_in <= 24'b010110100111011010011000;
#10000;
data_in <= 24'b010001010110000110000100;
#10000;
data_in <= 24'b010000000101011101111101;
#10000;
data_in <= 24'b010000100101011101111101;
#10000;
data_in <= 24'b010010100101100110000000;
#10000;
data_in <= 24'b010100110110000010000110;
#10000;
data_in <= 24'b011000000111110010011011;
#10000;
data_in <= 24'b011000110111111110100001;
#10000;
data_in <= 24'b010101000111001010010101;
#10000;
data_in <= 24'b010000100110000010000011;
#10000;
data_in <= 24'b010000000101101001111111;
#10000;
data_in <= 24'b010000110101101010000000;
#10000;
data_in <= 24'b010010100101101110000010;
#10000;
data_in <= 24'b010100010110000110000110;
#10000;
data_in <= 24'b011000010111110010011110;
#10000;
data_in <= 24'b010111100111110110011110;
#10000;
data_in <= 24'b010011010110110110010000;
#10000;
data_in <= 24'b001111100101111010000001;
#10000;
data_in <= 24'b010000010101110010000001;
#10000;
data_in <= 24'b010001010101110010000010;
#10000;
data_in <= 24'b010010010101110010000010;
#10000;
data_in <= 24'b010011100110000010000101;
#10000;
data_in <= 24'b011000100111111010100000;
#10000;
data_in <= 24'b010110100111101010011101;
#10000;
data_in <= 24'b010010010110100110001101;
#10000;
data_in <= 24'b001110110101101101111111;
#10000;
data_in <= 24'b010000000101101110000000;
#10000;
data_in <= 24'b010000110101110110000010;
#10000;
data_in <= 24'b010001110101101010000000;
#10000;
data_in <= 24'b010011000101111010000011;
#10000;
data_in <= 24'b011000101000000010100011;
#10000;
data_in <= 24'b010101110111101010011100;
#10000;
data_in <= 24'b010001000110011010001010;
#10000;
data_in <= 24'b001110000101100001111100;
#10000;
data_in <= 24'b001111010101101001111111;
#10000;
data_in <= 24'b010000100101110010000001;
#10000;
data_in <= 24'b010001100101100101111111;
#10000;
data_in <= 24'b010010100101110010000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010010100101011101110111;
#10000;
data_in <= 24'b010011010101100001110110;
#10000;
data_in <= 24'b010011100101100101110111;
#10000;
data_in <= 24'b010011100101110001111001;
#10000;
data_in <= 24'b010100000101111001111011;
#10000;
data_in <= 24'b010100010101111101111100;
#10000;
data_in <= 24'b010100010110000010000000;
#10000;
data_in <= 24'b010100100110000110000001;
#10000;
data_in <= 24'b010011110101101001111010;
#10000;
data_in <= 24'b010100000101101101111001;
#10000;
data_in <= 24'b010100010101110001111010;
#10000;
data_in <= 24'b010100010101111101111100;
#10000;
data_in <= 24'b010100100110000001111101;
#10000;
data_in <= 24'b010101000110001001111111;
#10000;
data_in <= 24'b010100110110001010000010;
#10000;
data_in <= 24'b010101010110010010000100;
#10000;
data_in <= 24'b010100000101110001111110;
#10000;
data_in <= 24'b010100010101111001111110;
#10000;
data_in <= 24'b010100110110000010000000;
#10000;
data_in <= 24'b010101000110000110000001;
#10000;
data_in <= 24'b010101010110001110000000;
#10000;
data_in <= 24'b010101000110010010000001;
#10000;
data_in <= 24'b010101110110011110000100;
#10000;
data_in <= 24'b010110010110100110000110;
#10000;
data_in <= 24'b010100000101111110000000;
#10000;
data_in <= 24'b010100100110000110000001;
#10000;
data_in <= 24'b010101100110001110000011;
#10000;
data_in <= 24'b010101000110001110000011;
#10000;
data_in <= 24'b010101000110010010000001;
#10000;
data_in <= 24'b010101100110011010000011;
#10000;
data_in <= 24'b010110010110100110000110;
#10000;
data_in <= 24'b010111000110110010001001;
#10000;
data_in <= 24'b010011100101111110000000;
#10000;
data_in <= 24'b010100010110001110000010;
#10000;
data_in <= 24'b010101010110010010000100;
#10000;
data_in <= 24'b010100110110010110000100;
#10000;
data_in <= 24'b010100100110010010000001;
#10000;
data_in <= 24'b010101000110011010000011;
#10000;
data_in <= 24'b010110010110101110001000;
#10000;
data_in <= 24'b010111100111000010001101;
#10000;
data_in <= 24'b010011000101111110000000;
#10000;
data_in <= 24'b010011110110001110000010;
#10000;
data_in <= 24'b010101000110011010000101;
#10000;
data_in <= 24'b010101000110011010000101;
#10000;
data_in <= 24'b010100110110010110000100;
#10000;
data_in <= 24'b010101100110100010000101;
#10000;
data_in <= 24'b010111000110111010001011;
#10000;
data_in <= 24'b011000010111010010001111;
#10000;
data_in <= 24'b010011000101111110000010;
#10000;
data_in <= 24'b010011110110010010000100;
#10000;
data_in <= 24'b010100110110011010000111;
#10000;
data_in <= 24'b010100110110011110000110;
#10000;
data_in <= 24'b010100100110011010000101;
#10000;
data_in <= 24'b010101010110101010000110;
#10000;
data_in <= 24'b010111010111001010001110;
#10000;
data_in <= 24'b011001000111100110010100;
#10000;
data_in <= 24'b010010110101111110000010;
#10000;
data_in <= 24'b010011110110010010000100;
#10000;
data_in <= 24'b010100110110100010001000;
#10000;
data_in <= 24'b010100110110100010001000;
#10000;
data_in <= 24'b010101000110100010000111;
#10000;
data_in <= 24'b010101110110101110001010;
#10000;
data_in <= 24'b010111110111010010010000;
#10000;
data_in <= 24'b011001110111110010010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000000111001010010001;
#10000;
data_in <= 24'b011100101000011010100101;
#10000;
data_in <= 24'b100010111001111010111111;
#10000;
data_in <= 24'b100111111011010011010100;
#10000;
data_in <= 24'b101011011100010011100100;
#10000;
data_in <= 24'b101101111100111111101101;
#10000;
data_in <= 24'b101110011101001011110010;
#10000;
data_in <= 24'b101110001101001011110000;
#10000;
data_in <= 24'b011000110111010110010100;
#10000;
data_in <= 24'b011101101000100010100111;
#10000;
data_in <= 24'b100011011010000111000000;
#10000;
data_in <= 24'b101000011011011011010101;
#10000;
data_in <= 24'b101100001100010111100101;
#10000;
data_in <= 24'b101110011101000111101111;
#10000;
data_in <= 24'b101111011101010011110100;
#10000;
data_in <= 24'b101111001101010011110010;
#10000;
data_in <= 24'b011001110111100110010110;
#10000;
data_in <= 24'b011110101000110010101001;
#10000;
data_in <= 24'b100100001010010111000001;
#10000;
data_in <= 24'b101001001011101011010110;
#10000;
data_in <= 24'b101100111100100011100111;
#10000;
data_in <= 24'b101111011101001111101111;
#10000;
data_in <= 24'b110000011101011011110101;
#10000;
data_in <= 24'b110000001101011011110010;
#10000;
data_in <= 24'b011010110111110110011010;
#10000;
data_in <= 24'b011111101001000010101101;
#10000;
data_in <= 24'b100100111010100011000100;
#10000;
data_in <= 24'b101001111011110011010111;
#10000;
data_in <= 24'b101101101100101111100110;
#10000;
data_in <= 24'b110000001101011111110001;
#10000;
data_in <= 24'b110001001101100111110100;
#10000;
data_in <= 24'b110001001101100111110100;
#10000;
data_in <= 24'b011100001000001110011110;
#10000;
data_in <= 24'b100000101001010110110000;
#10000;
data_in <= 24'b100110011010110011000111;
#10000;
data_in <= 24'b101011001100000011011001;
#10000;
data_in <= 24'b101110101100111011100111;
#10000;
data_in <= 24'b110000111101100111110010;
#10000;
data_in <= 24'b110010011101110111110110;
#10000;
data_in <= 24'b110010101101110011110011;
#10000;
data_in <= 24'b011101011000100010100011;
#10000;
data_in <= 24'b100001101001101010110011;
#10000;
data_in <= 24'b100111011011000111001010;
#10000;
data_in <= 24'b101011111100010011011010;
#10000;
data_in <= 24'b101111101101001111101001;
#10000;
data_in <= 24'b110010001101110111110011;
#10000;
data_in <= 24'b110011001110000111110111;
#10000;
data_in <= 24'b110011101110001011110100;
#10000;
data_in <= 24'b011110111000111010101001;
#10000;
data_in <= 24'b100011001010000010111001;
#10000;
data_in <= 24'b101000101011011011001111;
#10000;
data_in <= 24'b101101001100100111011111;
#10000;
data_in <= 24'b110000101101011111101101;
#10000;
data_in <= 24'b110011001110000111110110;
#10000;
data_in <= 24'b110100001110010111111010;
#10000;
data_in <= 24'b110100101110011011110111;
#10000;
data_in <= 24'b011111101001000110101100;
#10000;
data_in <= 24'b100011111010001110111100;
#10000;
data_in <= 24'b101001011011101011010000;
#10000;
data_in <= 24'b101101111100110011100010;
#10000;
data_in <= 24'b110001011101101011101111;
#10000;
data_in <= 24'b110011111110010011111001;
#10000;
data_in <= 24'b110100111110100111111011;
#10000;
data_in <= 24'b110101011110100111111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101100101100111011101100;
#10000;
data_in <= 24'b101100111100111111101101;
#10000;
data_in <= 24'b101100001100111011101011;
#10000;
data_in <= 24'b101011001100101011100111;
#10000;
data_in <= 24'b101010001100011111100110;
#10000;
data_in <= 24'b101010011100100011100111;
#10000;
data_in <= 24'b101001101100100011100110;
#10000;
data_in <= 24'b101001001100010111100110;
#10000;
data_in <= 24'b101110011101000111101111;
#10000;
data_in <= 24'b101110001101001111101110;
#10000;
data_in <= 24'b101101111101001011101101;
#10000;
data_in <= 24'b101100101100111111101010;
#10000;
data_in <= 24'b101101001101000111101100;
#10000;
data_in <= 24'b101110001101010011110010;
#10000;
data_in <= 24'b101110011101011111110100;
#10000;
data_in <= 24'b101101111101010111110010;
#10000;
data_in <= 24'b110000011101011011110001;
#10000;
data_in <= 24'b110000011101100011110010;
#10000;
data_in <= 24'b110000001101011111110001;
#10000;
data_in <= 24'b101111101101010111101111;
#10000;
data_in <= 24'b101111111101100011110010;
#10000;
data_in <= 24'b110001011101110111111001;
#10000;
data_in <= 24'b110001011110000011111011;
#10000;
data_in <= 24'b110000111101111011111001;
#10000;
data_in <= 24'b110010101101110011110011;
#10000;
data_in <= 24'b110010101101110011110011;
#10000;
data_in <= 24'b110010001101101011110001;
#10000;
data_in <= 24'b110001001101100011110001;
#10000;
data_in <= 24'b110001011101101111110100;
#10000;
data_in <= 24'b110010101101111111111010;
#10000;
data_in <= 24'b110010101110000111111011;
#10000;
data_in <= 24'b110001011101110111111001;
#10000;
data_in <= 24'b110011101101110111110000;
#10000;
data_in <= 24'b110011111101111011110001;
#10000;
data_in <= 24'b110011101101110111110000;
#10000;
data_in <= 24'b110011011101111011110011;
#10000;
data_in <= 24'b110011111110000111111000;
#10000;
data_in <= 24'b110101001110010111111111;
#10000;
data_in <= 24'b110100011110010011111111;
#10000;
data_in <= 24'b110010101101111111111011;
#10000;
data_in <= 24'b110011101101110011101110;
#10000;
data_in <= 24'b110100101101111111101111;
#10000;
data_in <= 24'b110100101110000011110010;
#10000;
data_in <= 24'b110101011110010011110111;
#10000;
data_in <= 24'b110110001110100111111110;
#10000;
data_in <= 24'b110110101110110011111111;
#10000;
data_in <= 24'b110101001110011111111111;
#10000;
data_in <= 24'b110010111110000011111100;
#10000;
data_in <= 24'b110100101110000111110001;
#10000;
data_in <= 24'b110101111110010011110010;
#10000;
data_in <= 24'b110101111110011011110110;
#10000;
data_in <= 24'b110101111110011111111000;
#10000;
data_in <= 24'b110110001110100111111110;
#10000;
data_in <= 24'b110101001110011011111101;
#10000;
data_in <= 24'b110001011101101011110101;
#10000;
data_in <= 24'b101110001100111011101010;
#10000;
data_in <= 24'b110110011110101011110111;
#10000;
data_in <= 24'b110110111110101111111000;
#10000;
data_in <= 24'b110110011110100111111001;
#10000;
data_in <= 24'b110101011110011111111000;
#10000;
data_in <= 24'b110011011110001011110111;
#10000;
data_in <= 24'b110000101101100111101111;
#10000;
data_in <= 24'b101011101100011011100010;
#10000;
data_in <= 24'b100111011011011111010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101000011100010011100101;
#10000;
data_in <= 24'b101001011100101111101011;
#10000;
data_in <= 24'b101001011100101111101101;
#10000;
data_in <= 24'b101000011100011111101001;
#10000;
data_in <= 24'b101000001100100011101011;
#10000;
data_in <= 24'b101001001100110011101111;
#10000;
data_in <= 24'b100111111100011111101010;
#10000;
data_in <= 24'b100101101011110111100011;
#10000;
data_in <= 24'b101101101101011011110011;
#10000;
data_in <= 24'b101100101101010011110001;
#10000;
data_in <= 24'b101011101101001011110000;
#10000;
data_in <= 24'b101011101101001011110000;
#10000;
data_in <= 24'b101011101101010011110100;
#10000;
data_in <= 24'b101010001100111111101111;
#10000;
data_in <= 24'b100101101011110111011101;
#10000;
data_in <= 24'b100001001010101011001101;
#10000;
data_in <= 24'b110000011101110111111011;
#10000;
data_in <= 24'b101110111101100111110110;
#10000;
data_in <= 24'b101101101101010111110100;
#10000;
data_in <= 24'b101101101101010111110110;
#10000;
data_in <= 24'b101010111100101111101110;
#10000;
data_in <= 24'b100101001011011111011001;
#10000;
data_in <= 24'b011110111001111011000000;
#10000;
data_in <= 24'b011010011000110110110001;
#10000;
data_in <= 24'b110000111101110111111011;
#10000;
data_in <= 24'b101111001101100011110111;
#10000;
data_in <= 24'b101101111101001011110100;
#10000;
data_in <= 24'b101011011100100111101100;
#10000;
data_in <= 24'b100100011010111111010010;
#10000;
data_in <= 24'b011011101000111010110010;
#10000;
data_in <= 24'b010111000111110010100000;
#10000;
data_in <= 24'b010110110111101010100001;
#10000;
data_in <= 24'b110010001101110111111100;
#10000;
data_in <= 24'b101110011101000011110000;
#10000;
data_in <= 24'b101010011100001011100100;
#10000;
data_in <= 24'b100101101011000011010100;
#10000;
data_in <= 24'b011110101001010010111001;
#10000;
data_in <= 24'b010110110111010110011101;
#10000;
data_in <= 24'b010100100110110010010100;
#10000;
data_in <= 24'b010101110111001110011100;
#10000;
data_in <= 24'b101111011101001011110010;
#10000;
data_in <= 24'b101001001011101011011101;
#10000;
data_in <= 24'b100010101010001011000110;
#10000;
data_in <= 24'b011110001001001010110111;
#10000;
data_in <= 24'b011010101000001110101011;
#10000;
data_in <= 24'b010110010111001110011011;
#10000;
data_in <= 24'b010100110110110010010110;
#10000;
data_in <= 24'b010101010111000010011100;
#10000;
data_in <= 24'b100110111011010011010100;
#10000;
data_in <= 24'b100001111010001011000100;
#10000;
data_in <= 24'b011100111000110110110010;
#10000;
data_in <= 24'b011001111000000110101001;
#10000;
data_in <= 24'b011000010111101110100011;
#10000;
data_in <= 24'b010110110111011110100000;
#10000;
data_in <= 24'b010110100111010110100001;
#10000;
data_in <= 24'b010110110111011010100010;
#10000;
data_in <= 24'b011111101001101010111100;
#10000;
data_in <= 24'b011101111001010110111000;
#10000;
data_in <= 24'b011011111000110010110011;
#10000;
data_in <= 24'b011001101000001110101010;
#10000;
data_in <= 24'b010111010111101110100100;
#10000;
data_in <= 24'b010110110111100110100010;
#10000;
data_in <= 24'b011000010111111010101010;
#10000;
data_in <= 24'b011001111000010010110000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100011111011001011011101;
#10000;
data_in <= 24'b011111101001111111001100;
#10000;
data_in <= 24'b011010011000101010110111;
#10000;
data_in <= 24'b010111000111110110101010;
#10000;
data_in <= 24'b010110100111101110101000;
#10000;
data_in <= 24'b011000011000001010101111;
#10000;
data_in <= 24'b011100001001001011000000;
#10000;
data_in <= 24'b011111111010001011001110;
#10000;
data_in <= 24'b011101101001100111000001;
#10000;
data_in <= 24'b011001011000011110110010;
#10000;
data_in <= 24'b010110000111101010100101;
#10000;
data_in <= 24'b010111010111111110101010;
#10000;
data_in <= 24'b011011001000110110111010;
#10000;
data_in <= 24'b011110011001101011000111;
#10000;
data_in <= 24'b011111111010000011001101;
#10000;
data_in <= 24'b100000101010001111010000;
#10000;
data_in <= 24'b011000011000000110101010;
#10000;
data_in <= 24'b010101100111011010100001;
#10000;
data_in <= 24'b010101000111010010011111;
#10000;
data_in <= 24'b011001101000011010110001;
#10000;
data_in <= 24'b011111111001111111001010;
#10000;
data_in <= 24'b100010101010101011010101;
#10000;
data_in <= 24'b100000111010001111001110;
#10000;
data_in <= 24'b011110001001100011000011;
#10000;
data_in <= 24'b010100100111001010011101;
#10000;
data_in <= 24'b010101000111010010011111;
#10000;
data_in <= 24'b010111010111110110101000;
#10000;
data_in <= 24'b011100001001000010111011;
#10000;
data_in <= 24'b100000001010000011001011;
#10000;
data_in <= 24'b100000101010001011001101;
#10000;
data_in <= 24'b011101111001010011000000;
#10000;
data_in <= 24'b011010101000011110110011;
#10000;
data_in <= 24'b010011100110101110010111;
#10000;
data_in <= 24'b010111000111100110100110;
#10000;
data_in <= 24'b011011101000101110110111;
#10000;
data_in <= 24'b011101111001010011000000;
#10000;
data_in <= 24'b011101011001001010111110;
#10000;
data_in <= 24'b011011111000110010111000;
#10000;
data_in <= 24'b011010101000011010101111;
#10000;
data_in <= 24'b011001011000000110101010;
#10000;
data_in <= 24'b010110100111010010100010;
#10000;
data_in <= 24'b011010011000011010110011;
#10000;
data_in <= 24'b011110001001010111000001;
#10000;
data_in <= 24'b011101111001001010111110;
#10000;
data_in <= 24'b011010011000010010110000;
#10000;
data_in <= 24'b011000000111100110100011;
#10000;
data_in <= 24'b010111100111011110100001;
#10000;
data_in <= 24'b010111110111100110100001;
#10000;
data_in <= 24'b011001111000000110101111;
#10000;
data_in <= 24'b011011111000100110110111;
#10000;
data_in <= 24'b011100111000111010111010;
#10000;
data_in <= 24'b011011111000100010110100;
#10000;
data_in <= 24'b011001010111111010101000;
#10000;
data_in <= 24'b011000010111101010100010;
#10000;
data_in <= 24'b011000010111011110100000;
#10000;
data_in <= 24'b010111110111011010011100;
#10000;
data_in <= 24'b011001101000000110101101;
#10000;
data_in <= 24'b011010001000000110101101;
#10000;
data_in <= 24'b011001010111111010101010;
#10000;
data_in <= 24'b011001010111110110100111;
#10000;
data_in <= 24'b011010101000001110101011;
#10000;
data_in <= 24'b011100011000100010101110;
#10000;
data_in <= 24'b011100011000011110101011;
#10000;
data_in <= 24'b011011000111111110100100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100000111010010011010001;
#10000;
data_in <= 24'b100000011010001011001111;
#10000;
data_in <= 24'b011111111010000011001101;
#10000;
data_in <= 24'b011111101010000011001011;
#10000;
data_in <= 24'b011111001001110011000111;
#10000;
data_in <= 24'b011100111001001110111110;
#10000;
data_in <= 24'b011001011000010110110000;
#10000;
data_in <= 24'b010110110111101110100110;
#10000;
data_in <= 24'b011110111001110011001001;
#10000;
data_in <= 24'b011110011001101011000111;
#10000;
data_in <= 24'b011101101001100011000011;
#10000;
data_in <= 24'b011101111001011111000010;
#10000;
data_in <= 24'b011101011001010110111110;
#10000;
data_in <= 24'b011100001001000010111001;
#10000;
data_in <= 24'b011001111000011110110000;
#10000;
data_in <= 24'b011000011000000110101100;
#10000;
data_in <= 24'b011100111001001110111110;
#10000;
data_in <= 24'b011100001001000010111011;
#10000;
data_in <= 24'b011011001000110010110111;
#10000;
data_in <= 24'b011011001000100110110101;
#10000;
data_in <= 24'b011011001000101010110011;
#10000;
data_in <= 24'b011010101000100010110001;
#10000;
data_in <= 24'b011001111000010110101110;
#10000;
data_in <= 24'b011000011000000110101100;
#10000;
data_in <= 24'b011010101000011110110011;
#10000;
data_in <= 24'b011001101000001110101111;
#10000;
data_in <= 24'b011000100111111110101011;
#10000;
data_in <= 24'b010111110111110110100110;
#10000;
data_in <= 24'b010111110111101110100100;
#10000;
data_in <= 24'b010111000111101010100011;
#10000;
data_in <= 24'b010111010111100110100010;
#10000;
data_in <= 24'b010110010111011110100000;
#10000;
data_in <= 24'b010111000111100010100001;
#10000;
data_in <= 24'b010110010111010110011110;
#10000;
data_in <= 24'b010101100111001010011011;
#10000;
data_in <= 24'b010100110111000010010111;
#10000;
data_in <= 24'b010100110110110110010101;
#10000;
data_in <= 24'b010100000110110110010100;
#10000;
data_in <= 24'b010100000110101010010010;
#10000;
data_in <= 24'b010011010110100110010010;
#10000;
data_in <= 24'b010101010110111010010110;
#10000;
data_in <= 24'b010101000110110110010101;
#10000;
data_in <= 24'b010100010110101010010010;
#10000;
data_in <= 24'b010011100110100010001101;
#10000;
data_in <= 24'b010010110110010010001100;
#10000;
data_in <= 24'b010010010110001010001010;
#10000;
data_in <= 24'b010010000110000110001001;
#10000;
data_in <= 24'b010001100110000010001000;
#10000;
data_in <= 24'b011000010111011010011100;
#10000;
data_in <= 24'b010111100111001110011001;
#10000;
data_in <= 24'b010110010110111010010100;
#10000;
data_in <= 24'b010100110110100110001101;
#10000;
data_in <= 24'b010010110110001010001000;
#10000;
data_in <= 24'b010010000101111110000101;
#10000;
data_in <= 24'b010010000101111110000101;
#10000;
data_in <= 24'b010001100101111110000111;
#10000;
data_in <= 24'b011100101000010110101000;
#10000;
data_in <= 24'b011011011000000010100011;
#10000;
data_in <= 24'b011001010111100010011011;
#10000;
data_in <= 24'b010110100110111010010001;
#10000;
data_in <= 24'b010100100110011010001001;
#10000;
data_in <= 24'b010011010110000110000100;
#10000;
data_in <= 24'b010011010110000010000101;
#10000;
data_in <= 24'b010010010110000010000110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010100010111001010100000;
#10000;
data_in <= 24'b010011100110111110011101;
#10000;
data_in <= 24'b010011000110101110011000;
#10000;
data_in <= 24'b010011010110101110010100;
#10000;
data_in <= 24'b010011110110110010010011;
#10000;
data_in <= 24'b010011000110011010001010;
#10000;
data_in <= 24'b001111000101010101110101;
#10000;
data_in <= 24'b001011110100011001100000;
#10000;
data_in <= 24'b010101010111010010100001;
#10000;
data_in <= 24'b010100000111000110011110;
#10000;
data_in <= 24'b010011010110110110011000;
#10000;
data_in <= 24'b010010110110101110010100;
#10000;
data_in <= 24'b010100010110110110010110;
#10000;
data_in <= 24'b010100000110101110010000;
#10000;
data_in <= 24'b010000110101111010000000;
#10000;
data_in <= 24'b001110010101000101101111;
#10000;
data_in <= 24'b010101100111010110100010;
#10000;
data_in <= 24'b010100100111000110011110;
#10000;
data_in <= 24'b010011010110110110011000;
#10000;
data_in <= 24'b010010110110101110010100;
#10000;
data_in <= 24'b010100100110111010010111;
#10000;
data_in <= 24'b010101010111000010010101;
#10000;
data_in <= 24'b010011100110100010001100;
#10000;
data_in <= 24'b010010000110000001111110;
#10000;
data_in <= 24'b010100010111000110011100;
#10000;
data_in <= 24'b010011110110111110011010;
#10000;
data_in <= 24'b010011000110110010010111;
#10000;
data_in <= 24'b010011000110101010010011;
#10000;
data_in <= 24'b010011110110111010010101;
#10000;
data_in <= 24'b010101000111000110010110;
#10000;
data_in <= 24'b010100100110110010010000;
#10000;
data_in <= 24'b010011010110011010000110;
#10000;
data_in <= 24'b010011000110100110010101;
#10000;
data_in <= 24'b010010110110101110010110;
#10000;
data_in <= 24'b010011010110101010010110;
#10000;
data_in <= 24'b010011000110101010010011;
#10000;
data_in <= 24'b010011110110111010010101;
#10000;
data_in <= 24'b010100110111000010010101;
#10000;
data_in <= 24'b010100100110111010010001;
#10000;
data_in <= 24'b010011010110100010001010;
#10000;
data_in <= 24'b010001110110010110001110;
#10000;
data_in <= 24'b010010010110100110010010;
#10000;
data_in <= 24'b010011010110101110010100;
#10000;
data_in <= 24'b010011100110110010010101;
#10000;
data_in <= 24'b010100000110111110010110;
#10000;
data_in <= 24'b010100110111001010011001;
#10000;
data_in <= 24'b010100110111000010010101;
#10000;
data_in <= 24'b010100000110110010001111;
#10000;
data_in <= 24'b010010010110011010001101;
#10000;
data_in <= 24'b010011000110101010010011;
#10000;
data_in <= 24'b010011110110110110010110;
#10000;
data_in <= 24'b010100000110111010010111;
#10000;
data_in <= 24'b010100010111000110011010;
#10000;
data_in <= 24'b010101110111011010011101;
#10000;
data_in <= 24'b010110010111100010011111;
#10000;
data_in <= 24'b010110010111011010011011;
#10000;
data_in <= 24'b010011100110100110001110;
#10000;
data_in <= 24'b010011100110110110010100;
#10000;
data_in <= 24'b010100010111000010010111;
#10000;
data_in <= 24'b010100100111000010011001;
#10000;
data_in <= 24'b010100110111001110011100;
#10000;
data_in <= 24'b010110100111101010100011;
#10000;
data_in <= 24'b010111100111111010100111;
#10000;
data_in <= 24'b011000000111111110100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000010110010000000110110;
#10000;
data_in <= 24'b000001110001100100101010;
#10000;
data_in <= 24'b000010000001100000100101;
#10000;
data_in <= 24'b000101000010000000101010;
#10000;
data_in <= 24'b000110110010011000101110;
#10000;
data_in <= 24'b000110000010000000100111;
#10000;
data_in <= 24'b000010100001001100010111;
#10000;
data_in <= 24'b000000000000100100001101;
#10000;
data_in <= 24'b000111110011010001001111;
#10000;
data_in <= 24'b000100010010010000111001;
#10000;
data_in <= 24'b000001000001010000100101;
#10000;
data_in <= 24'b000001100001010000100000;
#10000;
data_in <= 24'b000100010001110000100100;
#10000;
data_in <= 24'b000101010001111100100110;
#10000;
data_in <= 24'b000101010001111000100010;
#10000;
data_in <= 24'b000100100001101100011111;
#10000;
data_in <= 24'b001110000100111101101001;
#10000;
data_in <= 24'b001000000011010101001011;
#10000;
data_in <= 24'b000001110001100000101011;
#10000;
data_in <= 24'b000000000000111000011011;
#10000;
data_in <= 24'b000001110001001100011101;
#10000;
data_in <= 24'b000100100001110000100011;
#10000;
data_in <= 24'b000110100010001100100111;
#10000;
data_in <= 24'b000111010010011000101010;
#10000;
data_in <= 24'b010001010101101101110111;
#10000;
data_in <= 24'b001100000100010101011011;
#10000;
data_in <= 24'b000101110010100000111101;
#10000;
data_in <= 24'b000010000001011100100111;
#10000;
data_in <= 24'b000001100001001000011110;
#10000;
data_in <= 24'b000010100001010100011101;
#10000;
data_in <= 24'b000100000001101000100001;
#10000;
data_in <= 24'b000101110001111100100110;
#10000;
data_in <= 24'b010010000110000001111110;
#10000;
data_in <= 24'b001110100101000001101001;
#10000;
data_in <= 24'b001001110011100101010000;
#10000;
data_in <= 24'b000101100010011000110111;
#10000;
data_in <= 24'b000010000001010100100011;
#10000;
data_in <= 24'b000000100000111000011010;
#10000;
data_in <= 24'b000010000001000100011010;
#10000;
data_in <= 24'b000011110001100000100001;
#10000;
data_in <= 24'b010011000110010110000101;
#10000;
data_in <= 24'b010001100101110001111000;
#10000;
data_in <= 24'b001101110100101101100100;
#10000;
data_in <= 24'b001000110011010001001001;
#10000;
data_in <= 24'b000011110001110100101111;
#10000;
data_in <= 24'b000000100000111100011101;
#10000;
data_in <= 24'b000001110001000100011011;
#10000;
data_in <= 24'b000100000001100100100011;
#10000;
data_in <= 24'b010101100111000110010011;
#10000;
data_in <= 24'b010100100110101010001000;
#10000;
data_in <= 24'b010001100101101101110110;
#10000;
data_in <= 24'b001101000100011001011101;
#10000;
data_in <= 24'b000111010010110000111111;
#10000;
data_in <= 24'b000010010001100000101000;
#10000;
data_in <= 24'b000001100001000100011111;
#10000;
data_in <= 24'b000010110001010000100001;
#10000;
data_in <= 24'b010111100111101010011101;
#10000;
data_in <= 24'b010110000111001110010101;
#10000;
data_in <= 24'b010100000110100010000110;
#10000;
data_in <= 24'b010000000101011001101111;
#10000;
data_in <= 24'b001010010011110001010001;
#10000;
data_in <= 24'b000100010010000100110010;
#10000;
data_in <= 24'b000000110001000000100000;
#10000;
data_in <= 24'b000000010000110000011010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000000010000100100010000;
#10000;
data_in <= 24'b000001100001000000010111;
#10000;
data_in <= 24'b000010110001010100011100;
#10000;
data_in <= 24'b000011000001100000011110;
#10000;
data_in <= 24'b000100010001110100100001;
#10000;
data_in <= 24'b000101110010001100100111;
#10000;
data_in <= 24'b000110000010010100100111;
#10000;
data_in <= 24'b000101010010001000100100;
#10000;
data_in <= 24'b000001100001000000010111;
#10000;
data_in <= 24'b000001110001000100011000;
#10000;
data_in <= 24'b000001110001001100011001;
#10000;
data_in <= 24'b000010010001010100011011;
#10000;
data_in <= 24'b000100100001111000100010;
#10000;
data_in <= 24'b000110100010100100101100;
#10000;
data_in <= 24'b000111010010110000101111;
#10000;
data_in <= 24'b000110110010101000101100;
#10000;
data_in <= 24'b000100000001101000100001;
#10000;
data_in <= 24'b000011010001011000011111;
#10000;
data_in <= 24'b000010010001001100011010;
#10000;
data_in <= 24'b000010010001010100011011;
#10000;
data_in <= 24'b000100110001111100100101;
#10000;
data_in <= 24'b000111110010101100101111;
#10000;
data_in <= 24'b001001000011000000110100;
#10000;
data_in <= 24'b001001000011000100110011;
#10000;
data_in <= 24'b000110000010000100101010;
#10000;
data_in <= 24'b000101010001111000100111;
#10000;
data_in <= 24'b000100010001101000100011;
#10000;
data_in <= 24'b000100010001101100100010;
#10000;
data_in <= 24'b000101100010001000101000;
#10000;
data_in <= 24'b000111100010101000110000;
#10000;
data_in <= 24'b001001100011001000111000;
#10000;
data_in <= 24'b001010010011010100111001;
#10000;
data_in <= 24'b000110010010000000101001;
#10000;
data_in <= 24'b000110110010001000101011;
#10000;
data_in <= 24'b000110110010010000101101;
#10000;
data_in <= 24'b000110110010010000101101;
#10000;
data_in <= 24'b000110110010010000101101;
#10000;
data_in <= 24'b001000000010101000110001;
#10000;
data_in <= 24'b001010100011010000111011;
#10000;
data_in <= 24'b001100110011111001000010;
#10000;
data_in <= 24'b000100000001100100100011;
#10000;
data_in <= 24'b000101110001110100101000;
#10000;
data_in <= 24'b000110110010010000101110;
#10000;
data_in <= 24'b000111100010011100110000;
#10000;
data_in <= 24'b000111010010011000101111;
#10000;
data_in <= 24'b001000000010100100110010;
#10000;
data_in <= 24'b001011000011010100111110;
#10000;
data_in <= 24'b001110000100001001001001;
#10000;
data_in <= 24'b000010010001000100011110;
#10000;
data_in <= 24'b000011000001010000100001;
#10000;
data_in <= 24'b000100100001101000100111;
#10000;
data_in <= 24'b000101110010000000101010;
#10000;
data_in <= 24'b000110000010000100101011;
#10000;
data_in <= 24'b000110100010001100101100;
#10000;
data_in <= 24'b001001110010111000110111;
#10000;
data_in <= 24'b001101000011101101000100;
#10000;
data_in <= 24'b000001010000111000011100;
#10000;
data_in <= 24'b000001010000110100011010;
#10000;
data_in <= 24'b000010000001000000011101;
#10000;
data_in <= 24'b000011010001010100100010;
#10000;
data_in <= 24'b000100000001100000100101;
#10000;
data_in <= 24'b000100110001110000100110;
#10000;
data_in <= 24'b000111100010010000101111;
#10000;
data_in <= 24'b001010000010111100111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000110110010011100100111;
#10000;
data_in <= 24'b001000100010110000101100;
#10000;
data_in <= 24'b001000110010101100101010;
#10000;
data_in <= 24'b001000000010011000100101;
#10000;
data_in <= 24'b001000000010010100100011;
#10000;
data_in <= 24'b001001100010100100100111;
#10000;
data_in <= 24'b001010110010110000101010;
#10000;
data_in <= 24'b001010010010101000100110;
#10000;
data_in <= 24'b000101100010010000100011;
#10000;
data_in <= 24'b000110110010011100100111;
#10000;
data_in <= 24'b000111110010101000101000;
#10000;
data_in <= 24'b001000010010011100100110;
#10000;
data_in <= 24'b001000010010011000100100;
#10000;
data_in <= 24'b001001000010011100100101;
#10000;
data_in <= 24'b001010000010100100100111;
#10000;
data_in <= 24'b001010010010101000100110;
#10000;
data_in <= 24'b000110110010011100100111;
#10000;
data_in <= 24'b000110110010011100100111;
#10000;
data_in <= 24'b000111100010100100100111;
#10000;
data_in <= 24'b001001000010101000101001;
#10000;
data_in <= 24'b001001000010100100101000;
#10000;
data_in <= 24'b001001000010011100100101;
#10000;
data_in <= 24'b001001100010011100100101;
#10000;
data_in <= 24'b001010010010101000101000;
#10000;
data_in <= 24'b001001110011001100110101;
#10000;
data_in <= 24'b001000010010101100101011;
#10000;
data_in <= 24'b000111110010011100100111;
#10000;
data_in <= 24'b001000110010100100101000;
#10000;
data_in <= 24'b001001100010101100101010;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001001100010011000100110;
#10000;
data_in <= 24'b001010000010100100100111;
#10000;
data_in <= 24'b001100100011101100111111;
#10000;
data_in <= 24'b001001110011000000110011;
#10000;
data_in <= 24'b000111110010011000101001;
#10000;
data_in <= 24'b000111110010010000100101;
#10000;
data_in <= 24'b001000110010011100101000;
#10000;
data_in <= 24'b001001000010100000101001;
#10000;
data_in <= 24'b001001010010011100101000;
#10000;
data_in <= 24'b001001010010011100100111;
#10000;
data_in <= 24'b001111000100010001001011;
#10000;
data_in <= 24'b001101010011111001000010;
#10000;
data_in <= 24'b001010100011000000110101;
#10000;
data_in <= 24'b001000010010011000101001;
#10000;
data_in <= 24'b001000000010001100100111;
#10000;
data_in <= 24'b001000110010011000101010;
#10000;
data_in <= 24'b001001000010011100101011;
#10000;
data_in <= 24'b001000100010010100101001;
#10000;
data_in <= 24'b010011110101011001011111;
#10000;
data_in <= 24'b010100100101101001100001;
#10000;
data_in <= 24'b010010010100111101010110;
#10000;
data_in <= 24'b001100010011011100111100;
#10000;
data_in <= 24'b001001000010100000101101;
#10000;
data_in <= 24'b001001000010100000101101;
#10000;
data_in <= 24'b001001100010101000101111;
#10000;
data_in <= 24'b001000110010011100101100;
#10000;
data_in <= 24'b011001000110101001110101;
#10000;
data_in <= 24'b011011110111011001111111;
#10000;
data_in <= 24'b011010000110110101110110;
#10000;
data_in <= 24'b010001100100101101010100;
#10000;
data_in <= 24'b001010100010111100111000;
#10000;
data_in <= 24'b001001010010101100110010;
#10000;
data_in <= 24'b001001110010110000110101;
#10000;
data_in <= 24'b001000110010100100110000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010100100110000001110111;
#10000;
data_in <= 24'b001101100100010001011011;
#10000;
data_in <= 24'b000111100010101001000110;
#10000;
data_in <= 24'b000111100010101001000110;
#10000;
data_in <= 24'b001011100011101101011011;
#10000;
data_in <= 24'b010000100101000101110010;
#10000;
data_in <= 24'b010101010110100110001100;
#10000;
data_in <= 24'b011000010111101110011111;
#10000;
data_in <= 24'b010010010101011101101110;
#10000;
data_in <= 24'b001100000011111001010101;
#10000;
data_in <= 24'b000111000010100001000100;
#10000;
data_in <= 24'b000111010010101101001000;
#10000;
data_in <= 24'b001100000011110101011101;
#10000;
data_in <= 24'b010001000101010101110110;
#10000;
data_in <= 24'b010101110110110110010001;
#10000;
data_in <= 24'b011001000111111110100100;
#10000;
data_in <= 24'b001111010100110101100100;
#10000;
data_in <= 24'b001010010011100101010000;
#10000;
data_in <= 24'b000110100010100001000100;
#10000;
data_in <= 24'b000111110010110101001010;
#10000;
data_in <= 24'b001100010100000001100000;
#10000;
data_in <= 24'b010001100101100101111010;
#10000;
data_in <= 24'b010110100111000010010100;
#10000;
data_in <= 24'b011001101000000110100110;
#10000;
data_in <= 24'b001110010100100101100000;
#10000;
data_in <= 24'b001010000011101001010001;
#10000;
data_in <= 24'b000111110010111001001000;
#10000;
data_in <= 24'b001000110011001101010000;
#10000;
data_in <= 24'b001101000100011001100101;
#10000;
data_in <= 24'b010010000101110001111111;
#10000;
data_in <= 24'b010110010111000010010110;
#10000;
data_in <= 24'b011000111000000010100111;
#10000;
data_in <= 24'b001100110100011001011011;
#10000;
data_in <= 24'b001001110011110001010010;
#10000;
data_in <= 24'b001000100011001101001101;
#10000;
data_in <= 24'b001001100011100001010101;
#10000;
data_in <= 24'b001101100100100101101010;
#10000;
data_in <= 24'b010010010101111110000010;
#10000;
data_in <= 24'b010110100111010010011001;
#10000;
data_in <= 24'b011000111000001010101001;
#10000;
data_in <= 24'b001011010100001001010111;
#10000;
data_in <= 24'b001001110011110001010010;
#10000;
data_in <= 24'b001001000011100001010001;
#10000;
data_in <= 24'b001010000011110101011001;
#10000;
data_in <= 24'b001110000100110101101101;
#10000;
data_in <= 24'b010011000110001010000110;
#10000;
data_in <= 24'b010111000111011110011100;
#10000;
data_in <= 24'b011001001000001010101011;
#10000;
data_in <= 24'b001010110100001101010111;
#10000;
data_in <= 24'b001010000011111101010101;
#10000;
data_in <= 24'b001001100011110001010101;
#10000;
data_in <= 24'b001010100011111101011011;
#10000;
data_in <= 24'b001110000100110101101101;
#10000;
data_in <= 24'b010010010110000110000101;
#10000;
data_in <= 24'b010110100111010010011100;
#10000;
data_in <= 24'b011000010111111110101000;
#10000;
data_in <= 24'b001011100100010101011011;
#10000;
data_in <= 24'b001011000100001101011001;
#10000;
data_in <= 24'b001010010011111001011001;
#10000;
data_in <= 24'b001010100100000001011100;
#10000;
data_in <= 24'b001101000100101101101011;
#10000;
data_in <= 24'b010001010101110110000001;
#10000;
data_in <= 24'b010101010110111110010111;
#10000;
data_in <= 24'b010110110111100110100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010111100111101110100000;
#10000;
data_in <= 24'b010100000111001010010110;
#10000;
data_in <= 24'b010000100110001110001010;
#10000;
data_in <= 24'b001110010101101010000001;
#10000;
data_in <= 24'b001110110101100001111101;
#10000;
data_in <= 24'b010000000101101001111111;
#10000;
data_in <= 24'b010001110101101001111111;
#10000;
data_in <= 24'b010010000101101001111111;
#10000;
data_in <= 24'b010111100111111010100010;
#10000;
data_in <= 24'b010100000111000110011000;
#10000;
data_in <= 24'b010000000110010010001010;
#10000;
data_in <= 24'b001110000101100110000000;
#10000;
data_in <= 24'b001110100101011101111100;
#10000;
data_in <= 24'b010000100101100101111111;
#10000;
data_in <= 24'b010010000101101110000000;
#10000;
data_in <= 24'b010010010101101110000000;
#10000;
data_in <= 24'b010111110111111010100101;
#10000;
data_in <= 24'b010011110111001110011001;
#10000;
data_in <= 24'b001111110110001110001001;
#10000;
data_in <= 24'b001101110101100001111111;
#10000;
data_in <= 24'b001110110101011001111011;
#10000;
data_in <= 24'b010000010101100001111110;
#10000;
data_in <= 24'b010010010101101110000000;
#10000;
data_in <= 24'b010011000101110010000001;
#10000;
data_in <= 24'b010111110111111110101000;
#10000;
data_in <= 24'b010100000111001110011011;
#10000;
data_in <= 24'b001111110110001010001010;
#10000;
data_in <= 24'b001101100101011101111110;
#10000;
data_in <= 24'b001110010101010001111001;
#10000;
data_in <= 24'b010000100101011101111101;
#10000;
data_in <= 24'b010010110101101110000000;
#10000;
data_in <= 24'b010011110101110010000010;
#10000;
data_in <= 24'b010111101000000110101001;
#10000;
data_in <= 24'b010100000111010010011100;
#10000;
data_in <= 24'b001111110110001010001010;
#10000;
data_in <= 24'b001101110101011001111101;
#10000;
data_in <= 24'b001110100101010001111001;
#10000;
data_in <= 24'b010000110101011001111100;
#10000;
data_in <= 24'b010011010101101010000000;
#10000;
data_in <= 24'b010100010101110110000001;
#10000;
data_in <= 24'b010111101000000010101011;
#10000;
data_in <= 24'b010100000111001110011110;
#10000;
data_in <= 24'b001111110110001010001010;
#10000;
data_in <= 24'b001101110101011001111101;
#10000;
data_in <= 24'b001110100101001101111011;
#10000;
data_in <= 24'b010001000101011001111011;
#10000;
data_in <= 24'b010011100101100101111111;
#10000;
data_in <= 24'b010100000101110010000000;
#10000;
data_in <= 24'b010111101000000010101011;
#10000;
data_in <= 24'b010100000111001110011110;
#10000;
data_in <= 24'b010000000110001110001011;
#10000;
data_in <= 24'b001110000101011101111110;
#10000;
data_in <= 24'b001111010101001101111100;
#10000;
data_in <= 24'b010001000101011001111011;
#10000;
data_in <= 24'b010011100101100101111111;
#10000;
data_in <= 24'b010100010101101001111111;
#10000;
data_in <= 24'b011000001000000010101011;
#10000;
data_in <= 24'b010100010111010010011100;
#10000;
data_in <= 24'b010000100110001010001011;
#10000;
data_in <= 24'b001110010101100001111111;
#10000;
data_in <= 24'b001111010101010001111010;
#10000;
data_in <= 24'b010001010101011101111100;
#10000;
data_in <= 24'b010010110101100101111101;
#10000;
data_in <= 24'b010011110101101101111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010011010110000110000100;
#10000;
data_in <= 24'b010100010110010110001000;
#10000;
data_in <= 24'b010100010110011010000110;
#10000;
data_in <= 24'b010101000110100110001001;
#10000;
data_in <= 24'b010101100110101110001010;
#10000;
data_in <= 24'b010100110110100010000111;
#10000;
data_in <= 24'b010110100110111110001011;
#10000;
data_in <= 24'b011011011000001010011101;
#10000;
data_in <= 24'b010011010110000010000011;
#10000;
data_in <= 24'b010100010110010110001000;
#10000;
data_in <= 24'b010100010110011010000110;
#10000;
data_in <= 24'b010100110110100010001000;
#10000;
data_in <= 24'b010101100110101110001010;
#10000;
data_in <= 24'b010100110110100010000111;
#10000;
data_in <= 24'b010110110110111110001110;
#10000;
data_in <= 24'b011011111000010010100000;
#10000;
data_in <= 24'b010011010110000010000011;
#10000;
data_in <= 24'b010100010110010010000111;
#10000;
data_in <= 24'b010100100110010110000110;
#10000;
data_in <= 24'b010101000110011110001000;
#10000;
data_in <= 24'b010101100110100110001010;
#10000;
data_in <= 24'b010101000110100010000111;
#10000;
data_in <= 24'b010111010111001010010001;
#10000;
data_in <= 24'b011100101000100010100100;
#10000;
data_in <= 24'b010011100101111010000010;
#10000;
data_in <= 24'b010100010110010010000111;
#10000;
data_in <= 24'b010100100110010110000110;
#10000;
data_in <= 24'b010100110110011010000111;
#10000;
data_in <= 24'b010101100110100110001010;
#10000;
data_in <= 24'b010101100110100110001010;
#10000;
data_in <= 24'b011000010111011010010101;
#10000;
data_in <= 24'b011110001000110110101100;
#10000;
data_in <= 24'b010011100101111010000010;
#10000;
data_in <= 24'b010100110110001110000111;
#10000;
data_in <= 24'b010101000110010010001000;
#10000;
data_in <= 24'b010101010110010110001001;
#10000;
data_in <= 24'b010101110110101010001011;
#10000;
data_in <= 24'b010110010110110010001101;
#10000;
data_in <= 24'b011010000111101110011100;
#10000;
data_in <= 24'b100000011001010010110101;
#10000;
data_in <= 24'b010011110101110110000001;
#10000;
data_in <= 24'b010100100110001010000110;
#10000;
data_in <= 24'b010101000110010010001000;
#10000;
data_in <= 24'b010101100110011010001010;
#10000;
data_in <= 24'b010110100110101110001100;
#10000;
data_in <= 24'b010111000110111110010000;
#10000;
data_in <= 24'b011011111000001010100011;
#10000;
data_in <= 24'b100010101001110110111110;
#10000;
data_in <= 24'b010100000101110001111110;
#10000;
data_in <= 24'b010101000110001110000100;
#10000;
data_in <= 24'b010101100110010010001000;
#10000;
data_in <= 24'b010101110110011110001011;
#10000;
data_in <= 24'b010111000110110010010000;
#10000;
data_in <= 24'b011000100111001010010110;
#10000;
data_in <= 24'b011101001000011110101010;
#10000;
data_in <= 24'b100100101010010111001000;
#10000;
data_in <= 24'b010011100101110101111110;
#10000;
data_in <= 24'b010100100110010010000011;
#10000;
data_in <= 24'b010101000110010110000110;
#10000;
data_in <= 24'b010101110110100010001001;
#10000;
data_in <= 24'b010111010110110110010001;
#10000;
data_in <= 24'b011000100111010110011000;
#10000;
data_in <= 24'b011110001000101110101110;
#10000;
data_in <= 24'b100101011010100111001100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100000101001011110110010;
#10000;
data_in <= 24'b100101001010101011000011;
#10000;
data_in <= 24'b101010111100001011011000;
#10000;
data_in <= 24'b101110111101001011101000;
#10000;
data_in <= 24'b110010001101110111110010;
#10000;
data_in <= 24'b110100001110010111111010;
#10000;
data_in <= 24'b110100111110100011111101;
#10000;
data_in <= 24'b110100111110100111111011;
#10000;
data_in <= 24'b100001001001100110110101;
#10000;
data_in <= 24'b100101101010101111000110;
#10000;
data_in <= 24'b101011001100001011011011;
#10000;
data_in <= 24'b101111001101001111101001;
#10000;
data_in <= 24'b110001101101110111110011;
#10000;
data_in <= 24'b110011101110010111111011;
#10000;
data_in <= 24'b110101001110100111111111;
#10000;
data_in <= 24'b110101001110101011111100;
#10000;
data_in <= 24'b100011001010001010111110;
#10000;
data_in <= 24'b100111011011010011001110;
#10000;
data_in <= 24'b101100101100100111100011;
#10000;
data_in <= 24'b110000001101100011110000;
#10000;
data_in <= 24'b110010011110000111111001;
#10000;
data_in <= 24'b110100001110100011111111;
#10000;
data_in <= 24'b110100111110100111111111;
#10000;
data_in <= 24'b110100011110100111111111;
#10000;
data_in <= 24'b100101101010101111001010;
#10000;
data_in <= 24'b101001101011110011011000;
#10000;
data_in <= 24'b101110011100111111101011;
#10000;
data_in <= 24'b110001001101101011110110;
#10000;
data_in <= 24'b110010011101111111111011;
#10000;
data_in <= 24'b110010011110000111111101;
#10000;
data_in <= 24'b110010101110000111111011;
#10000;
data_in <= 24'b110001011101111011111000;
#10000;
data_in <= 24'b100111011011001011010010;
#10000;
data_in <= 24'b101011001100000111100000;
#10000;
data_in <= 24'b101110011101000111101111;
#10000;
data_in <= 24'b110000001101100011110110;
#10000;
data_in <= 24'b110000001101100011110110;
#10000;
data_in <= 24'b101111001101011011110100;
#10000;
data_in <= 24'b101110001101000011101110;
#10000;
data_in <= 24'b101100011100101111101001;
#10000;
data_in <= 24'b101001101011101111011011;
#10000;
data_in <= 24'b101011111100011011100110;
#10000;
data_in <= 24'b101110011100111111110010;
#10000;
data_in <= 24'b101110011101001011110010;
#10000;
data_in <= 24'b101101101100111111110001;
#10000;
data_in <= 24'b101100101100101111101101;
#10000;
data_in <= 24'b101011011100011011101000;
#10000;
data_in <= 24'b101001101100000111100011;
#10000;
data_in <= 24'b101010001011110011011111;
#10000;
data_in <= 24'b101011011100001111100110;
#10000;
data_in <= 24'b101100011100011111101011;
#10000;
data_in <= 24'b101011001100010111100111;
#10000;
data_in <= 24'b101010001100000011100100;
#10000;
data_in <= 24'b101001011011111111100011;
#10000;
data_in <= 24'b101001011011111111100011;
#10000;
data_in <= 24'b101001001011111011100010;
#10000;
data_in <= 24'b101000001011011011011010;
#10000;
data_in <= 24'b101000101011101011011110;
#10000;
data_in <= 24'b101000101011100111011111;
#10000;
data_in <= 24'b100110101011010011011001;
#10000;
data_in <= 24'b100101011011000011010101;
#10000;
data_in <= 24'b100110001011001111011000;
#10000;
data_in <= 24'b100110101011011111011110;
#10000;
data_in <= 24'b100111001011100111100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b110110011110110011111001;
#10000;
data_in <= 24'b110110001110101111111000;
#10000;
data_in <= 24'b110100111110100011110111;
#10000;
data_in <= 24'b110010101110001011110100;
#10000;
data_in <= 24'b110000101101110111110010;
#10000;
data_in <= 24'b101101101101001011101010;
#10000;
data_in <= 24'b101000011011111111011100;
#10000;
data_in <= 24'b100011111010111011001101;
#10000;
data_in <= 24'b110101101110110111111100;
#10000;
data_in <= 24'b110100011110101111111001;
#10000;
data_in <= 24'b110010001110001011110010;
#10000;
data_in <= 24'b101111101101100111101101;
#10000;
data_in <= 24'b101100101101000111101000;
#10000;
data_in <= 24'b101001011100011011100000;
#10000;
data_in <= 24'b100100101011010011010010;
#10000;
data_in <= 24'b011111111010010111000101;
#10000;
data_in <= 24'b110011101110100011111001;
#10000;
data_in <= 24'b110001111110001111110100;
#10000;
data_in <= 24'b101111001101101011101101;
#10000;
data_in <= 24'b101011101100111011100101;
#10000;
data_in <= 24'b101001001100010111011111;
#10000;
data_in <= 24'b100101111011101111011001;
#10000;
data_in <= 24'b100001111010110111001101;
#10000;
data_in <= 24'b011101111001111111000010;
#10000;
data_in <= 24'b101111111101101111110011;
#10000;
data_in <= 24'b101110001101011111101110;
#10000;
data_in <= 24'b101011111100111011100111;
#10000;
data_in <= 24'b101001011100011011100000;
#10000;
data_in <= 24'b100111101100000011011110;
#10000;
data_in <= 24'b100101001011100111011011;
#10000;
data_in <= 24'b100001111010110111010000;
#10000;
data_in <= 24'b011101111010000111000110;
#10000;
data_in <= 24'b101100001100101111100110;
#10000;
data_in <= 24'b101011011100101011100101;
#10000;
data_in <= 24'b101001111100010011100011;
#10000;
data_in <= 24'b100111111100000011100001;
#10000;
data_in <= 24'b100110111011111011100000;
#10000;
data_in <= 24'b100101001011100111011111;
#10000;
data_in <= 24'b100001111010111011010101;
#10000;
data_in <= 24'b011110011010000111001011;
#10000;
data_in <= 24'b101000111011111111011110;
#10000;
data_in <= 24'b101000111011111011100000;
#10000;
data_in <= 24'b101000001011110011011111;
#10000;
data_in <= 24'b100110111011101111011111;
#10000;
data_in <= 24'b100110011011101011100001;
#10000;
data_in <= 24'b100101011011011111100010;
#10000;
data_in <= 24'b100001111010110011011000;
#10000;
data_in <= 24'b011110101010000111001101;
#10000;
data_in <= 24'b100111001011011011011010;
#10000;
data_in <= 24'b100111001011011011011011;
#10000;
data_in <= 24'b100110101011010011011100;
#10000;
data_in <= 24'b100110011011010111011110;
#10000;
data_in <= 24'b100110101011011111100011;
#10000;
data_in <= 24'b100101111011100011100101;
#10000;
data_in <= 24'b100011101011000011011110;
#10000;
data_in <= 24'b100000101010011011010100;
#10000;
data_in <= 24'b100101111011001011010111;
#10000;
data_in <= 24'b100110001011001011010111;
#10000;
data_in <= 24'b100101111011000111011001;
#10000;
data_in <= 24'b100101111011001111011100;
#10000;
data_in <= 24'b100110111011100011100100;
#10000;
data_in <= 24'b100111011011110111101000;
#10000;
data_in <= 24'b100110001011100011100011;
#10000;
data_in <= 24'b100011101011000011011011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011111001001110010111111;
#10000;
data_in <= 24'b011101101001100010111100;
#10000;
data_in <= 24'b011011011000111010110101;
#10000;
data_in <= 24'b010111111000001010101010;
#10000;
data_in <= 24'b010101100111100110100001;
#10000;
data_in <= 24'b010101000111011110011111;
#10000;
data_in <= 24'b010110110111101110100100;
#10000;
data_in <= 24'b011000011000000110101010;
#10000;
data_in <= 24'b011101001001100010111100;
#10000;
data_in <= 24'b011011101001001110111001;
#10000;
data_in <= 24'b011001001000100010110000;
#10000;
data_in <= 24'b010110000111110010100100;
#10000;
data_in <= 24'b010011110111001110011011;
#10000;
data_in <= 24'b010011100111001010011010;
#10000;
data_in <= 24'b010100110111011010011110;
#10000;
data_in <= 24'b010110110111110010100011;
#10000;
data_in <= 24'b011011001001001110111001;
#10000;
data_in <= 24'b011001001000110110110100;
#10000;
data_in <= 24'b010110011000001010101001;
#10000;
data_in <= 24'b010100000111011110011110;
#10000;
data_in <= 24'b010010010111000010010110;
#10000;
data_in <= 24'b010010010111000010010110;
#10000;
data_in <= 24'b010011110111010010011010;
#10000;
data_in <= 24'b010101100111100010011100;
#10000;
data_in <= 24'b011010011001001010111001;
#10000;
data_in <= 24'b011000001000101110110010;
#10000;
data_in <= 24'b010101100111111110100110;
#10000;
data_in <= 24'b010011100111010110011100;
#10000;
data_in <= 24'b010010100111000110010111;
#10000;
data_in <= 24'b010011010111001110010110;
#10000;
data_in <= 24'b010100100111011010011010;
#10000;
data_in <= 24'b010110000111101110011101;
#10000;
data_in <= 24'b011010101001001010111100;
#10000;
data_in <= 24'b011000011000100110110011;
#10000;
data_in <= 24'b010101110111111010100101;
#10000;
data_in <= 24'b010011100111010110011011;
#10000;
data_in <= 24'b010011110111001110010111;
#10000;
data_in <= 24'b010101000111011110011001;
#10000;
data_in <= 24'b010110100111101110011100;
#10000;
data_in <= 24'b010111110111111010011111;
#10000;
data_in <= 24'b011100001001010111000001;
#10000;
data_in <= 24'b011001011000101010110110;
#10000;
data_in <= 24'b010101110111111010100101;
#10000;
data_in <= 24'b010100010111010110011011;
#10000;
data_in <= 24'b010100110111011010011000;
#10000;
data_in <= 24'b010110010111101010011011;
#10000;
data_in <= 24'b011000010111111010011101;
#10000;
data_in <= 24'b011000100111111110011110;
#10000;
data_in <= 24'b011110101001110011001010;
#10000;
data_in <= 24'b011011011001000010111100;
#10000;
data_in <= 24'b010111101000000110101001;
#10000;
data_in <= 24'b010101110111100110011101;
#10000;
data_in <= 24'b010110100111100110011010;
#10000;
data_in <= 24'b011000000111110110011100;
#10000;
data_in <= 24'b011001010111111110011101;
#10000;
data_in <= 24'b011001010111111110011101;
#10000;
data_in <= 24'b100000101010010011001111;
#10000;
data_in <= 24'b011101101001011010111111;
#10000;
data_in <= 24'b011001101000010110101100;
#10000;
data_in <= 24'b010111100111101110100000;
#10000;
data_in <= 24'b011000000111110010011111;
#10000;
data_in <= 24'b011000110111111010100000;
#10000;
data_in <= 24'b011001100111111110011111;
#10000;
data_in <= 24'b011001110111111010011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010111000111100010100001;
#10000;
data_in <= 24'b010111110111100010100010;
#10000;
data_in <= 24'b011001100111111010101000;
#10000;
data_in <= 24'b011100011000011110110000;
#10000;
data_in <= 24'b011110011000111110110011;
#10000;
data_in <= 24'b011111001001000010110011;
#10000;
data_in <= 24'b011111111001001010110011;
#10000;
data_in <= 24'b100000111001011010110111;
#10000;
data_in <= 24'b010110000111010010011101;
#10000;
data_in <= 24'b011000110111110010100100;
#10000;
data_in <= 24'b011100001000011010101111;
#10000;
data_in <= 24'b011111011001001110110111;
#10000;
data_in <= 24'b100001101001101010111101;
#10000;
data_in <= 24'b100010111001111010111111;
#10000;
data_in <= 24'b100011101010000010111111;
#10000;
data_in <= 24'b100011111001111110111100;
#10000;
data_in <= 24'b010110110111100010011111;
#10000;
data_in <= 24'b011001111000000110100110;
#10000;
data_in <= 24'b011100101000101010101110;
#10000;
data_in <= 24'b011111001001000010110011;
#10000;
data_in <= 24'b100001111001101010111011;
#10000;
data_in <= 24'b100101111010011111000100;
#10000;
data_in <= 24'b100111001010101011000110;
#10000;
data_in <= 24'b100110101010011111000001;
#10000;
data_in <= 24'b011000000111110010011111;
#10000;
data_in <= 24'b011010011000000110100101;
#10000;
data_in <= 24'b011011011000001110100110;
#10000;
data_in <= 24'b011100101000011110100110;
#10000;
data_in <= 24'b100001101001011010110011;
#10000;
data_in <= 24'b100111001010101111000101;
#10000;
data_in <= 24'b101000111010111111000111;
#10000;
data_in <= 24'b100111011010100010111100;
#10000;
data_in <= 24'b010111000111011110011001;
#10000;
data_in <= 24'b011001000111110110011111;
#10000;
data_in <= 24'b011011001000000110100000;
#10000;
data_in <= 24'b011100111000100010100100;
#10000;
data_in <= 24'b100010001001011110110001;
#10000;
data_in <= 24'b100101101010010010111010;
#10000;
data_in <= 24'b100011111001101010101110;
#10000;
data_in <= 24'b011111101000100010011001;
#10000;
data_in <= 24'b010111000111010110010101;
#10000;
data_in <= 24'b011001100111110110011101;
#10000;
data_in <= 24'b011011111000010010100011;
#10000;
data_in <= 24'b011101011000100010100011;
#10000;
data_in <= 24'b011110001000100010011111;
#10000;
data_in <= 24'b011011000111101010001101;
#10000;
data_in <= 24'b010100010101101101101100;
#10000;
data_in <= 24'b001101100011111101001101;
#10000;
data_in <= 24'b011000100111101110011011;
#10000;
data_in <= 24'b011001100111111010011100;
#10000;
data_in <= 24'b011010000111111010011010;
#10000;
data_in <= 24'b011000100111011010001111;
#10000;
data_in <= 24'b010100100110000001110110;
#10000;
data_in <= 24'b001101010100000101010011;
#10000;
data_in <= 24'b000101110010000000101110;
#10000;
data_in <= 24'b000000100000101100010101;
#10000;
data_in <= 24'b011010011000000110011111;
#10000;
data_in <= 24'b011001100111101110011010;
#10000;
data_in <= 24'b010111010111001010001101;
#10000;
data_in <= 24'b010011000101110101110111;
#10000;
data_in <= 24'b001100010011111101010101;
#10000;
data_in <= 24'b000100110001111100110001;
#10000;
data_in <= 24'b000000110000111000011100;
#10000;
data_in <= 24'b000000000000100000010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011110001000101010101001;
#10000;
data_in <= 24'b011100111000010110100100;
#10000;
data_in <= 24'b011010110111110110011100;
#10000;
data_in <= 24'b011000010111001110010010;
#10000;
data_in <= 24'b010110000110100110001010;
#10000;
data_in <= 24'b010100010110010010000101;
#10000;
data_in <= 24'b010011110110001010000101;
#10000;
data_in <= 24'b010011010110000110000100;
#10000;
data_in <= 24'b100001011001001110101111;
#10000;
data_in <= 24'b011101111000010110100001;
#10000;
data_in <= 24'b011001100111010010010000;
#10000;
data_in <= 24'b010110100110100010000100;
#10000;
data_in <= 24'b010011110101111101111100;
#10000;
data_in <= 24'b010010000101100001110101;
#10000;
data_in <= 24'b010001010101010001110100;
#10000;
data_in <= 24'b010000110101011001110111;
#10000;
data_in <= 24'b100010011001010110101101;
#10000;
data_in <= 24'b011011010111101010010000;
#10000;
data_in <= 24'b010100000101110001110100;
#10000;
data_in <= 24'b010000100100111001100110;
#10000;
data_in <= 24'b001101100100001101011101;
#10000;
data_in <= 24'b001010010011100001010010;
#10000;
data_in <= 24'b001001110011010101010001;
#10000;
data_in <= 24'b001010000011101001010111;
#10000;
data_in <= 24'b011101011000000010010100;
#10000;
data_in <= 24'b010100110101110101101111;
#10000;
data_in <= 24'b001100010011101001001110;
#10000;
data_in <= 24'b001000010010110001000000;
#10000;
data_in <= 24'b000101110010010000111010;
#10000;
data_in <= 24'b000010100001100000101110;
#10000;
data_in <= 24'b000010010001011100101110;
#10000;
data_in <= 24'b000010110001111000111001;
#10000;
data_in <= 24'b010001110100111101100000;
#10000;
data_in <= 24'b001010010011001001000000;
#10000;
data_in <= 24'b000100000001100000101001;
#10000;
data_in <= 24'b000010010001001100100100;
#10000;
data_in <= 24'b000010010001001100100101;
#10000;
data_in <= 24'b000000100000110100100001;
#10000;
data_in <= 24'b000001000001000100100111;
#10000;
data_in <= 24'b000010100001110000110011;
#10000;
data_in <= 24'b000100010001100100100110;
#10000;
data_in <= 24'b000000110000101100011000;
#10000;
data_in <= 24'b000000000000010100010010;
#10000;
data_in <= 24'b000000110000110000011010;
#10000;
data_in <= 24'b000010110001001100100100;
#10000;
data_in <= 24'b000011100001100000101010;
#10000;
data_in <= 24'b000101010010000100110011;
#10000;
data_in <= 24'b000111000010110101000010;
#10000;
data_in <= 24'b000000000000010000001110;
#10000;
data_in <= 24'b000000000000011000010001;
#10000;
data_in <= 24'b000010100001000000011011;
#10000;
data_in <= 24'b000101100001111100101001;
#10000;
data_in <= 24'b000111110010100000110101;
#10000;
data_in <= 24'b001001000010111100111101;
#10000;
data_in <= 24'b001011000011100101001001;
#10000;
data_in <= 24'b001011110100000001010011;
#10000;
data_in <= 24'b000000100000101100011000;
#10000;
data_in <= 24'b000100000001100100100110;
#10000;
data_in <= 24'b001000100010101100111000;
#10000;
data_in <= 24'b001011010011100001000110;
#10000;
data_in <= 24'b001100110100000001010000;
#10000;
data_in <= 24'b001101100100010001010110;
#10000;
data_in <= 24'b001110110100101001011101;
#10000;
data_in <= 24'b001111000100111001100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010100000110110010001111;
#10000;
data_in <= 24'b010011110110110010010001;
#10000;
data_in <= 24'b010100100111000110011000;
#10000;
data_in <= 24'b010110110111101010100001;
#10000;
data_in <= 24'b011000011000000110101010;
#10000;
data_in <= 24'b011000101000010110101101;
#10000;
data_in <= 24'b011000011000010010101100;
#10000;
data_in <= 24'b011000101000001010101011;
#10000;
data_in <= 24'b001101110101001001110100;
#10000;
data_in <= 24'b010000000101111010000001;
#10000;
data_in <= 24'b010011110110111110010011;
#10000;
data_in <= 24'b010111100111111110100110;
#10000;
data_in <= 24'b011001111000101010110010;
#10000;
data_in <= 24'b011010111000110110111000;
#10000;
data_in <= 24'b011011001000111010111001;
#10000;
data_in <= 24'b011011001000111010111001;
#10000;
data_in <= 24'b001000000011100101011001;
#10000;
data_in <= 24'b001101000101001001110101;
#10000;
data_in <= 24'b010100110111001110010111;
#10000;
data_in <= 24'b011010011000101010110001;
#10000;
data_in <= 24'b011100101001010110111101;
#10000;
data_in <= 24'b011100101001010111000000;
#10000;
data_in <= 24'b011100111001011011000010;
#10000;
data_in <= 24'b011100111001011011000010;
#10000;
data_in <= 24'b000110010011001101010001;
#10000;
data_in <= 24'b001110100101011001111000;
#10000;
data_in <= 24'b011001001000001010100101;
#10000;
data_in <= 24'b011110101001101111000010;
#10000;
data_in <= 24'b011111111010001011001010;
#10000;
data_in <= 24'b011110111001111011001010;
#10000;
data_in <= 24'b011101101001101011001000;
#10000;
data_in <= 24'b011101011001100111000111;
#10000;
data_in <= 24'b000111100011011001010010;
#10000;
data_in <= 24'b010000100101111101111110;
#10000;
data_in <= 24'b011011111000110110110000;
#10000;
data_in <= 24'b100001101010100011001100;
#10000;
data_in <= 24'b100010001010101111010011;
#10000;
data_in <= 24'b100000111010011011010010;
#10000;
data_in <= 24'b011111011010000111001111;
#10000;
data_in <= 24'b011110101001111011001100;
#10000;
data_in <= 24'b001000110011110001010110;
#10000;
data_in <= 24'b010001010110001010000001;
#10000;
data_in <= 24'b011100001000111110110000;
#10000;
data_in <= 24'b100001001010011011001010;
#10000;
data_in <= 24'b100010001010101111010011;
#10000;
data_in <= 24'b100000111010100011010100;
#10000;
data_in <= 24'b011111101010010111010010;
#10000;
data_in <= 24'b011110011001111111001111;
#10000;
data_in <= 24'b001110100101001101101101;
#10000;
data_in <= 24'b010101100111001110010010;
#10000;
data_in <= 24'b011110001001011110111000;
#10000;
data_in <= 24'b100001101010100011001100;
#10000;
data_in <= 24'b100010011010110111010101;
#10000;
data_in <= 24'b100010001010110111011001;
#10000;
data_in <= 24'b100000101010100011011000;
#10000;
data_in <= 24'b011110101010001011010010;
#10000;
data_in <= 24'b010111000111001010001110;
#10000;
data_in <= 24'b011100011000110110101100;
#10000;
data_in <= 24'b100011001010100011001010;
#10000;
data_in <= 24'b100101001011010011011000;
#10000;
data_in <= 24'b100101001011011111011111;
#10000;
data_in <= 24'b100100011011011011100010;
#10000;
data_in <= 24'b100010101011000011100000;
#10000;
data_in <= 24'b100000101010011111011001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000101000000110101000;
#10000;
data_in <= 24'b010111100111101010011101;
#10000;
data_in <= 24'b010110000111000110010001;
#10000;
data_in <= 24'b010100000110011010000010;
#10000;
data_in <= 24'b001110100100111001100111;
#10000;
data_in <= 24'b000111000010110101000010;
#10000;
data_in <= 24'b000001100001010000100110;
#10000;
data_in <= 24'b000000000000101100011011;
#10000;
data_in <= 24'b011010001000100010110001;
#10000;
data_in <= 24'b011000011000000010100111;
#10000;
data_in <= 24'b010110110111010110011001;
#10000;
data_in <= 24'b010101000110110010001010;
#10000;
data_in <= 24'b010001000101100101110100;
#10000;
data_in <= 24'b001011000011111001010101;
#10000;
data_in <= 24'b000100110010000100110111;
#10000;
data_in <= 24'b000000110001000100100011;
#10000;
data_in <= 24'b011011111001000110111100;
#10000;
data_in <= 24'b011010011000100110110010;
#10000;
data_in <= 24'b011001000111111110100100;
#10000;
data_in <= 24'b010111000111010110010111;
#10000;
data_in <= 24'b010101000110100110001000;
#10000;
data_in <= 24'b010000100101011001101111;
#10000;
data_in <= 24'b001001110011011101001110;
#10000;
data_in <= 24'b000100000001111100110010;
#10000;
data_in <= 24'b011100101001010111000001;
#10000;
data_in <= 24'b011100001001001010111101;
#10000;
data_in <= 24'b011011001000100110110000;
#10000;
data_in <= 24'b011001000111111010100010;
#10000;
data_in <= 24'b010111100111010110010101;
#10000;
data_in <= 24'b010100100110011110000011;
#10000;
data_in <= 24'b001110010100101001100100;
#10000;
data_in <= 24'b001000000011000101000110;
#10000;
data_in <= 24'b011100011001010111000011;
#10000;
data_in <= 24'b011100111001011011000010;
#10000;
data_in <= 24'b011100101001000010111001;
#10000;
data_in <= 24'b011010101000010110101010;
#10000;
data_in <= 24'b011000110111110010011110;
#10000;
data_in <= 24'b010110100110111110001110;
#10000;
data_in <= 24'b010001100101100101110100;
#10000;
data_in <= 24'b001100110100001101011010;
#10000;
data_in <= 24'b011101001001100011001000;
#10000;
data_in <= 24'b011101011001100011000100;
#10000;
data_in <= 24'b011100101001001010111101;
#10000;
data_in <= 24'b011011011000101010110001;
#10000;
data_in <= 24'b011001110111111110100011;
#10000;
data_in <= 24'b010111100111001110010010;
#10000;
data_in <= 24'b010011110110000101111110;
#10000;
data_in <= 24'b010000110101010001101110;
#10000;
data_in <= 24'b011110001001111011001110;
#10000;
data_in <= 24'b011100111001011111000101;
#10000;
data_in <= 24'b011011111001000010111101;
#10000;
data_in <= 24'b011011011000110010110011;
#10000;
data_in <= 24'b011010101000010010101000;
#10000;
data_in <= 24'b010111110111011010010110;
#10000;
data_in <= 24'b010101000110100010000111;
#10000;
data_in <= 24'b010011110110001101111100;
#10000;
data_in <= 24'b011111101010010011010100;
#10000;
data_in <= 24'b011100111001011111000111;
#10000;
data_in <= 24'b011011011000111010111100;
#10000;
data_in <= 24'b011011101000101110110111;
#10000;
data_in <= 24'b011011001000011010101110;
#10000;
data_in <= 24'b011000000111100010011100;
#10000;
data_in <= 24'b010110000110110010001111;
#10000;
data_in <= 24'b010101000110100110000101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000000100000101100011001;
#10000;
data_in <= 24'b000000110000110000011010;
#10000;
data_in <= 24'b000001010000111000011100;
#10000;
data_in <= 24'b000001100000111100011101;
#10000;
data_in <= 24'b000001010000110000011011;
#10000;
data_in <= 24'b000001100000111000011011;
#10000;
data_in <= 24'b000011010001010100100010;
#10000;
data_in <= 24'b000101010001111000101000;
#10000;
data_in <= 24'b000010000001001000100011;
#10000;
data_in <= 24'b000010010001010000100010;
#10000;
data_in <= 24'b000010100001010100100011;
#10000;
data_in <= 24'b000010110001010000100010;
#10000;
data_in <= 24'b000001110001000000011110;
#10000;
data_in <= 24'b000010100001000100100000;
#10000;
data_in <= 24'b000101000001101100101010;
#10000;
data_in <= 24'b001000000010100000110101;
#10000;
data_in <= 24'b000100010001111100110001;
#10000;
data_in <= 24'b000101000010000100110001;
#10000;
data_in <= 24'b000101010010001000110010;
#10000;
data_in <= 24'b000100110001110100101110;
#10000;
data_in <= 24'b000010110001010100100110;
#10000;
data_in <= 24'b000010110001001100100100;
#10000;
data_in <= 24'b000101110001111100110000;
#10000;
data_in <= 24'b001001010010111000111100;
#10000;
data_in <= 24'b000101000010010000110101;
#10000;
data_in <= 24'b000101100010010100110101;
#10000;
data_in <= 24'b000110010010100000111000;
#10000;
data_in <= 24'b000110000010010100110101;
#10000;
data_in <= 24'b000011010001101000101010;
#10000;
data_in <= 24'b000001110001000100100010;
#10000;
data_in <= 24'b000011010001011100101000;
#10000;
data_in <= 24'b000110110010010100110110;
#10000;
data_in <= 24'b000100010010001000110101;
#10000;
data_in <= 24'b000100110010001100110100;
#10000;
data_in <= 24'b000101110010011100111000;
#10000;
data_in <= 24'b000110100010100000111010;
#10000;
data_in <= 24'b000100000001111000110000;
#10000;
data_in <= 24'b000001100001001000100100;
#10000;
data_in <= 24'b000001100001001000100100;
#10000;
data_in <= 24'b000011100001101000101100;
#10000;
data_in <= 24'b000111010011000101000011;
#10000;
data_in <= 24'b000110100010110000111101;
#10000;
data_in <= 24'b000110110010110100111110;
#10000;
data_in <= 24'b001000100011001001000011;
#10000;
data_in <= 24'b000111010010110100111110;
#10000;
data_in <= 24'b000100100010000000110010;
#10000;
data_in <= 24'b000011110001101100101101;
#10000;
data_in <= 24'b000100110001111100110001;
#10000;
data_in <= 24'b001101100100110001011110;
#10000;
data_in <= 24'b001010000011110001001101;
#10000;
data_in <= 24'b000111110011001101000100;
#10000;
data_in <= 24'b001001010011011101001000;
#10000;
data_in <= 24'b001001110011011001001001;
#10000;
data_in <= 24'b000111010010110000111111;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
data_in <= 24'b000110010010011100111010;
#10000;
data_in <= 24'b010001110101110001110010;
#10000;
data_in <= 24'b001011110100010101010111;
#10000;
data_in <= 24'b000111100011000101000110;
#10000;
data_in <= 24'b000111110011001001000111;
#10000;
data_in <= 24'b001000000011001001001001;
#10000;
data_in <= 24'b000110000010101001000001;
#10000;
data_in <= 24'b000100010010001100111010;
#10000;
data_in <= 24'b000100100010010000111011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010011110101010101100010;
#10000;
data_in <= 24'b011110101000000010001011;
#10000;
data_in <= 24'b100011011001001110011110;
#10000;
data_in <= 24'b011100110111100110000100;
#10000;
data_in <= 24'b010011110101010101100000;
#10000;
data_in <= 24'b001101000011101101000100;
#10000;
data_in <= 24'b001001100010110000110111;
#10000;
data_in <= 24'b001001010010110000110101;
#10000;
data_in <= 24'b010110110110001001110001;
#10000;
data_in <= 24'b100000101000101010010111;
#10000;
data_in <= 24'b100101101001110110101100;
#10000;
data_in <= 24'b100010001001000010011101;
#10000;
data_in <= 24'b011011110111011110000100;
#10000;
data_in <= 24'b010100010101101001100111;
#10000;
data_in <= 24'b001100100011101101001000;
#10000;
data_in <= 24'b001000000010100100110110;
#10000;
data_in <= 24'b010011010101010101100110;
#10000;
data_in <= 24'b011100000111100110000111;
#10000;
data_in <= 24'b100010011001000110100010;
#10000;
data_in <= 24'b100011001001011110100101;
#10000;
data_in <= 24'b100010011001010010100010;
#10000;
data_in <= 24'b011101011000000010001110;
#10000;
data_in <= 24'b010011000101100101100111;
#10000;
data_in <= 24'b001011110011110001001010;
#10000;
data_in <= 24'b001100110011101101001100;
#10000;
data_in <= 24'b010101000101111001101111;
#10000;
data_in <= 24'b011100100111110010001101;
#10000;
data_in <= 24'b100000101000111110011111;
#10000;
data_in <= 24'b100011111001110010101100;
#10000;
data_in <= 24'b100001011001010010100100;
#10000;
data_in <= 24'b011010000111011010001000;
#10000;
data_in <= 24'b010011110101111101101111;
#10000;
data_in <= 24'b001001100011000001000010;
#10000;
data_in <= 24'b010010110101011101101001;
#10000;
data_in <= 24'b011011100111101010001100;
#10000;
data_in <= 24'b011111111000110110011111;
#10000;
data_in <= 24'b100010011001100110101010;
#10000;
data_in <= 24'b100000011001001110100100;
#10000;
data_in <= 24'b011011111000000010010011;
#10000;
data_in <= 24'b011000100111010010000101;
#10000;
data_in <= 24'b000110110010011100111001;
#10000;
data_in <= 24'b010001000101001001100100;
#10000;
data_in <= 24'b011010100111100010001010;
#10000;
data_in <= 24'b011110011000100110011010;
#10000;
data_in <= 24'b011110111000110010011111;
#10000;
data_in <= 24'b011100001000010010010110;
#10000;
data_in <= 24'b011000110111011110001001;
#10000;
data_in <= 24'b010111000111001010000100;
#10000;
data_in <= 24'b000100100010000000110011;
#10000;
data_in <= 24'b001110000100011001011001;
#10000;
data_in <= 24'b010110000110011101111010;
#10000;
data_in <= 24'b011000100111001110000110;
#10000;
data_in <= 24'b011000010111010010001001;
#10000;
data_in <= 24'b010101110110110010000001;
#10000;
data_in <= 24'b010011010110001001110111;
#10000;
data_in <= 24'b010010110110001101110111;
#10000;
data_in <= 24'b000100100010010000111011;
#10000;
data_in <= 24'b001100000100001101011000;
#10000;
data_in <= 24'b010001100101100101101110;
#10000;
data_in <= 24'b010011000101111101110100;
#10000;
data_in <= 24'b010011010110000001110101;
#10000;
data_in <= 24'b010001100101101001101100;
#10000;
data_in <= 24'b001111110101001101100101;
#10000;
data_in <= 24'b010000000101010001100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001100000100010001011101;
#10000;
data_in <= 24'b001010000011111001010111;
#10000;
data_in <= 24'b001001000011100101010100;
#10000;
data_in <= 24'b001001110011110001011011;
#10000;
data_in <= 24'b001011000100010101100111;
#10000;
data_in <= 24'b001110010101001101110111;
#10000;
data_in <= 24'b010011100110101110010010;
#10000;
data_in <= 24'b010111110111111010100101;
#10000;
data_in <= 24'b001100110100011101100000;
#10000;
data_in <= 24'b001010010011111101011000;
#10000;
data_in <= 24'b001000110011100001010100;
#10000;
data_in <= 24'b001000010011100101010111;
#10000;
data_in <= 24'b001010000100000101100011;
#10000;
data_in <= 24'b001101010101000101110100;
#10000;
data_in <= 24'b010010110110100010001101;
#10000;
data_in <= 24'b010111010111110010100011;
#10000;
data_in <= 24'b001101100100101001100011;
#10000;
data_in <= 24'b001011000100001001011011;
#10000;
data_in <= 24'b001000110011100001010100;
#10000;
data_in <= 24'b000111100011011001010100;
#10000;
data_in <= 24'b001000110011110001011100;
#10000;
data_in <= 24'b001100110100111101110010;
#10000;
data_in <= 24'b010010110110100010001101;
#10000;
data_in <= 24'b010111010111110010100011;
#10000;
data_in <= 24'b001101110100101101100100;
#10000;
data_in <= 24'b001011010100001101011100;
#10000;
data_in <= 24'b001000100011011101010010;
#10000;
data_in <= 24'b000110110011001101010001;
#10000;
data_in <= 24'b001000010011101001011010;
#10000;
data_in <= 24'b001100110100111101110010;
#10000;
data_in <= 24'b010011100110101110010000;
#10000;
data_in <= 24'b011000000111111110100110;
#10000;
data_in <= 24'b001100110100100001011110;
#10000;
data_in <= 24'b001010100100000001011001;
#10000;
data_in <= 24'b000111110011010001001111;
#10000;
data_in <= 24'b000101100010111001001100;
#10000;
data_in <= 24'b000111100011011101010111;
#10000;
data_in <= 24'b001100110100111101110010;
#10000;
data_in <= 24'b010011110110110010010001;
#10000;
data_in <= 24'b011001001000000110101000;
#10000;
data_in <= 24'b001011010100001001011000;
#10000;
data_in <= 24'b001010000011110001010101;
#10000;
data_in <= 24'b000111000011000101001100;
#10000;
data_in <= 24'b000101000010110001001010;
#10000;
data_in <= 24'b000111000011010101010101;
#10000;
data_in <= 24'b001101000100111001110010;
#10000;
data_in <= 24'b010100100110110110010010;
#10000;
data_in <= 24'b011000111000000010100111;
#10000;
data_in <= 24'b001011100100000001010111;
#10000;
data_in <= 24'b001010010011110101010110;
#10000;
data_in <= 24'b000111100011001101001110;
#10000;
data_in <= 24'b000110000010111001001010;
#10000;
data_in <= 24'b001000000011011101010111;
#10000;
data_in <= 24'b001101110101000101110101;
#10000;
data_in <= 24'b010100110110111010010011;
#10000;
data_in <= 24'b011000100111111110100100;
#10000;
data_in <= 24'b001100010100001101011010;
#10000;
data_in <= 24'b001011000100000101010111;
#10000;
data_in <= 24'b001001000011100001010001;
#10000;
data_in <= 24'b000111000011001001001110;
#10000;
data_in <= 24'b001000110011101001011010;
#10000;
data_in <= 24'b001110100101010101110111;
#10000;
data_in <= 24'b010101010111000110010100;
#10000;
data_in <= 24'b011000111000000010100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000111000000110101010;
#10000;
data_in <= 24'b010100000111000010011001;
#10000;
data_in <= 24'b001111110101110110000110;
#10000;
data_in <= 24'b001110100101011101111110;
#10000;
data_in <= 24'b001111000101011001111011;
#10000;
data_in <= 24'b010000100101100001111100;
#10000;
data_in <= 24'b010001110101101101111110;
#10000;
data_in <= 24'b010011000101111110000000;
#10000;
data_in <= 24'b011000101000000010101001;
#10000;
data_in <= 24'b010100100111000010011001;
#10000;
data_in <= 24'b010000110110000010000111;
#10000;
data_in <= 24'b001111010101100001111101;
#10000;
data_in <= 24'b001111000101011001111011;
#10000;
data_in <= 24'b001111110101011101111011;
#10000;
data_in <= 24'b010001010101101101111110;
#10000;
data_in <= 24'b010010110110001010000010;
#10000;
data_in <= 24'b010111110111110110100110;
#10000;
data_in <= 24'b010100100111000010011001;
#10000;
data_in <= 24'b010001010110001010001001;
#10000;
data_in <= 24'b001111100101100101111110;
#10000;
data_in <= 24'b001110110101010101111010;
#10000;
data_in <= 24'b001111100101011001111010;
#10000;
data_in <= 24'b010001100101110001111111;
#10000;
data_in <= 24'b010011100110001110000011;
#10000;
data_in <= 24'b010111010111101110100100;
#10000;
data_in <= 24'b010100110111000110011010;
#10000;
data_in <= 24'b010010000110010110001100;
#10000;
data_in <= 24'b001111110101101001111111;
#10000;
data_in <= 24'b001110110101010101111010;
#10000;
data_in <= 24'b001111100101011001111010;
#10000;
data_in <= 24'b010010010101110110000000;
#10000;
data_in <= 24'b010011110110010010000100;
#10000;
data_in <= 24'b010111000111101010100011;
#10000;
data_in <= 24'b010101000111001010011011;
#10000;
data_in <= 24'b010010010110011010001101;
#10000;
data_in <= 24'b001111110101101001111111;
#10000;
data_in <= 24'b001110110101010101111010;
#10000;
data_in <= 24'b001111110101011101111011;
#10000;
data_in <= 24'b010010010101110110000000;
#10000;
data_in <= 24'b010011100110001110000011;
#10000;
data_in <= 24'b010111100111110010100101;
#10000;
data_in <= 24'b010110000111010110011100;
#10000;
data_in <= 24'b010011000110011010001110;
#10000;
data_in <= 24'b010000000101101001111111;
#10000;
data_in <= 24'b001111010101010101111001;
#10000;
data_in <= 24'b010000110101100101111100;
#10000;
data_in <= 24'b010010010101111001111110;
#10000;
data_in <= 24'b010010100101111101111111;
#10000;
data_in <= 24'b011000100111111110100110;
#10000;
data_in <= 24'b010110010111011010011101;
#10000;
data_in <= 24'b010010110110010110001101;
#10000;
data_in <= 24'b001111110101100101111110;
#10000;
data_in <= 24'b001111100101011001111010;
#10000;
data_in <= 24'b010001010101101101111110;
#10000;
data_in <= 24'b010010010101111001111110;
#10000;
data_in <= 24'b010001110101110001111100;
#10000;
data_in <= 24'b011000111000000010100111;
#10000;
data_in <= 24'b010110100111011110011110;
#10000;
data_in <= 24'b010010110110011010001011;
#10000;
data_in <= 24'b001111110101100101111101;
#10000;
data_in <= 24'b001111110101011101111011;
#10000;
data_in <= 24'b010001100101110001111111;
#10000;
data_in <= 24'b010010010101111001111110;
#10000;
data_in <= 24'b010001100101100101111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010010110101111101111110;
#10000;
data_in <= 24'b010100000110010110000001;
#10000;
data_in <= 24'b010101010110100110001000;
#10000;
data_in <= 24'b010101010110100110001000;
#10000;
data_in <= 24'b010101110110101010001011;
#10000;
data_in <= 24'b011001000111100010011011;
#10000;
data_in <= 24'b011110111000111110110010;
#10000;
data_in <= 24'b100011101010000111000110;
#10000;
data_in <= 24'b010011100110010010000000;
#10000;
data_in <= 24'b010011110110011010000000;
#10000;
data_in <= 24'b010100010110011110000011;
#10000;
data_in <= 24'b010101010110101110000111;
#10000;
data_in <= 24'b010111000111000110010001;
#10000;
data_in <= 24'b011001100111101110011011;
#10000;
data_in <= 24'b011100001000001110101000;
#10000;
data_in <= 24'b011101101000100110101110;
#10000;
data_in <= 24'b010011110110010010000011;
#10000;
data_in <= 24'b010100100110100010000100;
#10000;
data_in <= 24'b010101100110101110000111;
#10000;
data_in <= 24'b010110000110110110001001;
#10000;
data_in <= 24'b010110010110110010001101;
#10000;
data_in <= 24'b010110100110110110001110;
#10000;
data_in <= 24'b010110100110110110010010;
#10000;
data_in <= 24'b010111000110111110010100;
#10000;
data_in <= 24'b010100010110011010000101;
#10000;
data_in <= 24'b010110000110111010001010;
#10000;
data_in <= 24'b010111000111000110001101;
#10000;
data_in <= 24'b010100110110011110000110;
#10000;
data_in <= 24'b010001010101100001111001;
#10000;
data_in <= 24'b001111100101000101110010;
#10000;
data_in <= 24'b010001000101011101111010;
#10000;
data_in <= 24'b010011000101111110000100;
#10000;
data_in <= 24'b010110000110110010001011;
#10000;
data_in <= 24'b010110000110110010001011;
#10000;
data_in <= 24'b010100110110010110000100;
#10000;
data_in <= 24'b010001000101011001110101;
#10000;
data_in <= 24'b001101000100010101100110;
#10000;
data_in <= 24'b001011110100000001100001;
#10000;
data_in <= 24'b001110000100100001101100;
#10000;
data_in <= 24'b010000000101001101110110;
#10000;
data_in <= 24'b010101110110101110001010;
#10000;
data_in <= 24'b010010100101111001111101;
#10000;
data_in <= 24'b001111000100111001101101;
#10000;
data_in <= 24'b001100000100001001100001;
#10000;
data_in <= 24'b001011100011111101100000;
#10000;
data_in <= 24'b001100100100001101100100;
#10000;
data_in <= 24'b001101100100011101101000;
#10000;
data_in <= 24'b001110010100100101101101;
#10000;
data_in <= 24'b010000110101011001110111;
#10000;
data_in <= 24'b001110100100101101101100;
#10000;
data_in <= 24'b001011110011111001011110;
#10000;
data_in <= 24'b001011000011101101011011;
#10000;
data_in <= 24'b001100110100001001100010;
#10000;
data_in <= 24'b001110110100101001101010;
#10000;
data_in <= 24'b001111100100110101101101;
#10000;
data_in <= 24'b001110110100110001101101;
#10000;
data_in <= 24'b001011010011111001011111;
#10000;
data_in <= 24'b001011000011111001011101;
#10000;
data_in <= 24'b001011100011110101011101;
#10000;
data_in <= 24'b001100000011111101011111;
#10000;
data_in <= 24'b001101010100010001100100;
#10000;
data_in <= 24'b001111000100110001101001;
#10000;
data_in <= 24'b010001010101001001110010;
#10000;
data_in <= 24'b010001100101010101110101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100100001010010111001011;
#10000;
data_in <= 24'b100001111001111011000100;
#10000;
data_in <= 24'b011111101001100011000000;
#10000;
data_in <= 24'b011111011001101011000001;
#10000;
data_in <= 24'b100000001001111111000110;
#10000;
data_in <= 24'b100001011010010011001011;
#10000;
data_in <= 24'b100010011010100111010010;
#10000;
data_in <= 24'b100011101010111011010111;
#10000;
data_in <= 24'b011100001000010110101011;
#10000;
data_in <= 24'b011010011000001110101000;
#10000;
data_in <= 24'b011010011000001110101011;
#10000;
data_in <= 24'b011011101000101010110011;
#10000;
data_in <= 24'b011100111001000110111010;
#10000;
data_in <= 24'b011101011001010110111110;
#10000;
data_in <= 24'b011110011001101111000110;
#10000;
data_in <= 24'b011111101010000111001001;
#10000;
data_in <= 24'b010101110110110010010010;
#10000;
data_in <= 24'b010110000110111110010101;
#10000;
data_in <= 24'b010111010111011010011110;
#10000;
data_in <= 24'b011001001000000110101000;
#10000;
data_in <= 24'b011010001000011010101111;
#10000;
data_in <= 24'b011010001000100010110001;
#10000;
data_in <= 24'b011010011000101110110110;
#10000;
data_in <= 24'b011011101001000110111001;
#10000;
data_in <= 24'b010100110110011010001100;
#10000;
data_in <= 24'b010101010110101010010000;
#10000;
data_in <= 24'b010110000111000110011001;
#10000;
data_in <= 24'b010111100111100010100000;
#10000;
data_in <= 24'b010111100111101010100011;
#10000;
data_in <= 24'b010110100111100010100001;
#10000;
data_in <= 24'b010110010111100110100100;
#10000;
data_in <= 24'b010111010111110110100110;
#10000;
data_in <= 24'b010011010110000010000101;
#10000;
data_in <= 24'b010011010110001010001000;
#10000;
data_in <= 24'b010011100110010010001101;
#10000;
data_in <= 24'b010011110110100010010000;
#10000;
data_in <= 24'b010011010110011010010000;
#10000;
data_in <= 24'b010010000110010010001101;
#10000;
data_in <= 24'b010001110110010010010000;
#10000;
data_in <= 24'b010010110110100110010010;
#10000;
data_in <= 24'b010001110101101001111101;
#10000;
data_in <= 24'b010001000101011101111100;
#10000;
data_in <= 24'b010000110101100001111110;
#10000;
data_in <= 24'b010001000101101010000011;
#10000;
data_in <= 24'b010000110101110010000100;
#10000;
data_in <= 24'b010000100101101110000101;
#10000;
data_in <= 24'b010001000101111110001011;
#10000;
data_in <= 24'b010010010110010110001110;
#10000;
data_in <= 24'b010001100101011001111010;
#10000;
data_in <= 24'b010000010101001101111000;
#10000;
data_in <= 24'b010000000101001101111000;
#10000;
data_in <= 24'b010001000101100101111111;
#10000;
data_in <= 24'b010010010101111110001000;
#10000;
data_in <= 24'b010011000110010110001101;
#10000;
data_in <= 24'b010100100110101010010100;
#10000;
data_in <= 24'b010101100111000010011000;
#10000;
data_in <= 24'b010010000101011101111000;
#10000;
data_in <= 24'b010000100101001001110110;
#10000;
data_in <= 24'b010000010101010001110111;
#10000;
data_in <= 24'b010010000101101110000000;
#10000;
data_in <= 24'b010100010110011010001100;
#10000;
data_in <= 24'b010101110110110110010110;
#10000;
data_in <= 24'b010111010111001110011100;
#10000;
data_in <= 24'b011000000111100110100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100010101010100111010000;
#10000;
data_in <= 24'b100011001010100111001110;
#10000;
data_in <= 24'b100011111010110011010001;
#10000;
data_in <= 24'b100101101011011011011010;
#10000;
data_in <= 24'b101001011100001111100110;
#10000;
data_in <= 24'b101011001100101011101101;
#10000;
data_in <= 24'b101010001100011011101001;
#10000;
data_in <= 24'b100111111011110111100000;
#10000;
data_in <= 24'b100000001001111111000110;
#10000;
data_in <= 24'b100001101010011011001010;
#10000;
data_in <= 24'b100011101010111011010001;
#10000;
data_in <= 24'b100110001011100111011010;
#10000;
data_in <= 24'b101010001100011111101000;
#10000;
data_in <= 24'b101101001101001111110010;
#10000;
data_in <= 24'b101101111101010111110010;
#10000;
data_in <= 24'b101100011100111111101100;
#10000;
data_in <= 24'b011100111001001010111001;
#10000;
data_in <= 24'b100000111010000011000101;
#10000;
data_in <= 24'b100100011010111111010010;
#10000;
data_in <= 24'b100110101011100111011010;
#10000;
data_in <= 24'b101001111100011011100111;
#10000;
data_in <= 24'b101110001101011111110110;
#10000;
data_in <= 24'b110000001101111111111110;
#10000;
data_in <= 24'b101111101101110111111100;
#10000;
data_in <= 24'b011010101000011110101110;
#10000;
data_in <= 24'b011111001001100110111110;
#10000;
data_in <= 24'b100011011010101111001110;
#10000;
data_in <= 24'b100101011011001111010110;
#10000;
data_in <= 24'b101000011100000011100001;
#10000;
data_in <= 24'b101100111101001011110001;
#10000;
data_in <= 24'b110000001101111111111110;
#10000;
data_in <= 24'b110000001110001011111111;
#10000;
data_in <= 24'b010111110111110010100001;
#10000;
data_in <= 24'b011100011000110110110000;
#10000;
data_in <= 24'b100000001001111011000001;
#10000;
data_in <= 24'b100010111010100111001100;
#10000;
data_in <= 24'b100101011011011011010111;
#10000;
data_in <= 24'b101001101100011111101000;
#10000;
data_in <= 24'b101101011101011011110111;
#10000;
data_in <= 24'b101110101101110111111110;
#10000;
data_in <= 24'b010110010111010010011001;
#10000;
data_in <= 24'b011000100111111010100001;
#10000;
data_in <= 24'b011100011000110110110000;
#10000;
data_in <= 24'b100000011001111111000010;
#10000;
data_in <= 24'b100011101010111111010000;
#10000;
data_in <= 24'b100111001011110111011110;
#10000;
data_in <= 24'b101010011100110011101101;
#10000;
data_in <= 24'b101100111101100111111001;
#10000;
data_in <= 24'b010110110111010110011010;
#10000;
data_in <= 24'b010110010111010110011000;
#10000;
data_in <= 24'b011001011000000110100100;
#10000;
data_in <= 24'b011111001001101010111101;
#10000;
data_in <= 24'b100011001010110011001111;
#10000;
data_in <= 24'b100101011011010111011000;
#10000;
data_in <= 24'b101000001100001111100101;
#10000;
data_in <= 24'b101011011101001011110100;
#10000;
data_in <= 24'b011000110111101010100000;
#10000;
data_in <= 24'b010110000111001010010110;
#10000;
data_in <= 24'b011000010111101110011111;
#10000;
data_in <= 24'b011111011001100110111100;
#10000;
data_in <= 24'b100011001010110011001111;
#10000;
data_in <= 24'b100011111011001011010100;
#10000;
data_in <= 24'b100101111011110011011110;
#10000;
data_in <= 24'b101001111100110111101111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100101001011001011010101;
#10000;
data_in <= 24'b100001011010000111000100;
#10000;
data_in <= 24'b011011111000101110101110;
#10000;
data_in <= 24'b011000000111101110100000;
#10000;
data_in <= 24'b010111110111100110011110;
#10000;
data_in <= 24'b011001010111111110100100;
#10000;
data_in <= 24'b011011101000100010101101;
#10000;
data_in <= 24'b011101111000110110110001;
#10000;
data_in <= 24'b100111001011100111011000;
#10000;
data_in <= 24'b100011011010101011001001;
#10000;
data_in <= 24'b011110101001010010111000;
#10000;
data_in <= 24'b011010111000011110101010;
#10000;
data_in <= 24'b011010101000001110101011;
#10000;
data_in <= 24'b011100011000101110110011;
#10000;
data_in <= 24'b011111011001010110111111;
#10000;
data_in <= 24'b100001101001110111000011;
#10000;
data_in <= 24'b101000101100000111100000;
#10000;
data_in <= 24'b100101101011010111010100;
#10000;
data_in <= 24'b100001111010001111000110;
#10000;
data_in <= 24'b011101111001010110111000;
#10000;
data_in <= 24'b011101101001000010111000;
#10000;
data_in <= 24'b011111011001101011000001;
#10000;
data_in <= 24'b100011011010011011010000;
#10000;
data_in <= 24'b100101111011000111010110;
#10000;
data_in <= 24'b101010001100101011101000;
#10000;
data_in <= 24'b100111101011111111100000;
#10000;
data_in <= 24'b100011111010111111010010;
#10000;
data_in <= 24'b100000011010000111000100;
#10000;
data_in <= 24'b011111011001110011000011;
#10000;
data_in <= 24'b100000111010001011001001;
#10000;
data_in <= 24'b100100001010111011010111;
#10000;
data_in <= 24'b100111011011101011100001;
#10000;
data_in <= 24'b101011101101000111110010;
#10000;
data_in <= 24'b101001101100100111101010;
#10000;
data_in <= 24'b100101111011101011011100;
#10000;
data_in <= 24'b100010101010110111001111;
#10000;
data_in <= 24'b100000101010011011001100;
#10000;
data_in <= 24'b100001011010100111001111;
#10000;
data_in <= 24'b100011101011000111011001;
#10000;
data_in <= 24'b100101111011100011011111;
#10000;
data_in <= 24'b101100101101100011111000;
#10000;
data_in <= 24'b101010011100111111110001;
#10000;
data_in <= 24'b100111001100001011100100;
#10000;
data_in <= 24'b100100011011011111011010;
#10000;
data_in <= 24'b100010101010111111010101;
#10000;
data_in <= 24'b100010001010111111010101;
#10000;
data_in <= 24'b100011011011000111011001;
#10000;
data_in <= 24'b100100001011010111011011;
#10000;
data_in <= 24'b101100001101011011111000;
#10000;
data_in <= 24'b101001111100111111110010;
#10000;
data_in <= 24'b100111001100010011100111;
#10000;
data_in <= 24'b100101001011110011011111;
#10000;
data_in <= 24'b100100001011011111011101;
#10000;
data_in <= 24'b100011001011011011011011;
#10000;
data_in <= 24'b100011001011001111011001;
#10000;
data_in <= 24'b100010111011001011011000;
#10000;
data_in <= 24'b101010111101001111110110;
#10000;
data_in <= 24'b101000101100110011101111;
#10000;
data_in <= 24'b100110011100001111100110;
#10000;
data_in <= 24'b100101001011111011100001;
#10000;
data_in <= 24'b100100101011110011100001;
#10000;
data_in <= 24'b100011111011100111011110;
#10000;
data_in <= 24'b100010111011010111011010;
#10000;
data_in <= 24'b100001101011000011010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011101111000101110101010;
#10000;
data_in <= 24'b011100111000010010011111;
#10000;
data_in <= 24'b010011010101101101110111;
#10000;
data_in <= 24'b001001000011001101001101;
#10000;
data_in <= 24'b000111010010101001000000;
#10000;
data_in <= 24'b000111010010101100111110;
#10000;
data_in <= 24'b000111110010101100111101;
#10000;
data_in <= 24'b001010000011010001000110;
#10000;
data_in <= 24'b100010001001110010111011;
#10000;
data_in <= 24'b010110100110101110000110;
#10000;
data_in <= 24'b001010010011011101010011;
#10000;
data_in <= 24'b000111110010111001001000;
#10000;
data_in <= 24'b001101000100001001011001;
#10000;
data_in <= 24'b010000000100111001100100;
#10000;
data_in <= 24'b010011000101101001110000;
#10000;
data_in <= 24'b010111000110101010000000;
#10000;
data_in <= 24'b100101001010100111001001;
#10000;
data_in <= 24'b010100100110011110000011;
#10000;
data_in <= 24'b001011110100000101011110;
#10000;
data_in <= 24'b010001110101101001110101;
#10000;
data_in <= 24'b011000000111000110001011;
#10000;
data_in <= 24'b011000000111001010001001;
#10000;
data_in <= 24'b011001010111010110001100;
#10000;
data_in <= 24'b011011101000000010010111;
#10000;
data_in <= 24'b100110011011010011010110;
#10000;
data_in <= 24'b011100101000101010101000;
#10000;
data_in <= 24'b011011001000010010100010;
#10000;
data_in <= 24'b100001111001110110111001;
#10000;
data_in <= 24'b100001101001110110110111;
#10000;
data_in <= 24'b011101011000101010100101;
#10000;
data_in <= 24'b011011111000010110011110;
#10000;
data_in <= 24'b011011101000010010011101;
#10000;
data_in <= 24'b100110111011100111011100;
#10000;
data_in <= 24'b100100011010111011001101;
#10000;
data_in <= 24'b100101111011010011010011;
#10000;
data_in <= 24'b100111001011100011010111;
#10000;
data_in <= 24'b100011101010101011001000;
#10000;
data_in <= 24'b100010111010011011000001;
#10000;
data_in <= 24'b100100001010101111000110;
#10000;
data_in <= 24'b100011101010011011000010;
#10000;
data_in <= 24'b100011011011000111010101;
#10000;
data_in <= 24'b100100111011011011011000;
#10000;
data_in <= 24'b100110011011100111011100;
#10000;
data_in <= 24'b100100111011010011010101;
#10000;
data_in <= 24'b100100101011000111010000;
#10000;
data_in <= 24'b100111001011101111011010;
#10000;
data_in <= 24'b101001111100010011100011;
#10000;
data_in <= 24'b101000101011111111011110;
#10000;
data_in <= 24'b100001111010111011010100;
#10000;
data_in <= 24'b100011001011010011010111;
#10000;
data_in <= 24'b100011101011010011010111;
#10000;
data_in <= 24'b100100001011011011011001;
#10000;
data_in <= 24'b100110101011111111100001;
#10000;
data_in <= 24'b100111111100001011100100;
#10000;
data_in <= 24'b101000001100000111100010;
#10000;
data_in <= 24'b101000111100010011100101;
#10000;
data_in <= 24'b100100001011101011011111;
#10000;
data_in <= 24'b100011101011100011011101;
#10000;
data_in <= 24'b100010101011001111011010;
#10000;
data_in <= 24'b100101101011110111100011;
#10000;
data_in <= 24'b101000101100100111101111;
#10000;
data_in <= 24'b100110101100000011100011;
#10000;
data_in <= 24'b100110001011110011100000;
#10000;
data_in <= 24'b101011011101001011110100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010000110100111101100001;
#10000;
data_in <= 24'b010000000100111001100001;
#10000;
data_in <= 24'b010000110101001001100101;
#10000;
data_in <= 24'b010001100101011101101100;
#10000;
data_in <= 24'b010001000101011001101101;
#10000;
data_in <= 24'b010001100101101001110011;
#10000;
data_in <= 24'b010101110110110010000111;
#10000;
data_in <= 24'b011010111000000110011101;
#10000;
data_in <= 24'b010111000110101010000000;
#10000;
data_in <= 24'b010100110110001101111010;
#10000;
data_in <= 24'b010011110110001101111100;
#10000;
data_in <= 24'b010101000110100110000100;
#10000;
data_in <= 24'b010111010111001110001111;
#10000;
data_in <= 24'b011001110111111110011101;
#10000;
data_in <= 24'b011110101001001110110011;
#10000;
data_in <= 24'b100011011010011011000110;
#10000;
data_in <= 24'b011000100111010010001011;
#10000;
data_in <= 24'b010110100110111010000111;
#10000;
data_in <= 24'b010111000111000010001001;
#10000;
data_in <= 24'b011010111000000010011011;
#10000;
data_in <= 24'b100000001001011010110010;
#10000;
data_in <= 24'b100100011010100111000111;
#10000;
data_in <= 24'b101000101011101111011011;
#10000;
data_in <= 24'b101100001100100111101001;
#10000;
data_in <= 24'b011010111000000010011011;
#10000;
data_in <= 24'b011010111000000010011011;
#10000;
data_in <= 24'b011101001000101110100101;
#10000;
data_in <= 24'b100010011001111110111011;
#10000;
data_in <= 24'b100111011011010111010011;
#10000;
data_in <= 24'b101010101100010011100010;
#10000;
data_in <= 24'b101100011100110111101100;
#10000;
data_in <= 24'b101110001101010011110011;
#10000;
data_in <= 24'b100100001010100011000100;
#10000;
data_in <= 24'b100101001010110011001000;
#10000;
data_in <= 24'b100111011011010111010001;
#10000;
data_in <= 24'b101010001100001011100000;
#10000;
data_in <= 24'b101100011100101111101001;
#10000;
data_in <= 24'b101100111100111111101110;
#10000;
data_in <= 24'b101101011101000011110010;
#10000;
data_in <= 24'b101101101101001011110001;
#10000;
data_in <= 24'b101010001100010011100011;
#10000;
data_in <= 24'b101010011100010111100011;
#10000;
data_in <= 24'b101011011100100111101000;
#10000;
data_in <= 24'b101100001100110011101011;
#10000;
data_in <= 24'b101100101100111011101101;
#10000;
data_in <= 24'b101100111101000011101111;
#10000;
data_in <= 24'b101101101101001011110100;
#10000;
data_in <= 24'b101110001101010011110110;
#10000;
data_in <= 24'b101010101100100111101010;
#10000;
data_in <= 24'b101010101100100111101000;
#10000;
data_in <= 24'b101011001100100011101010;
#10000;
data_in <= 24'b101011011100100111101011;
#10000;
data_in <= 24'b101100001100110011101110;
#10000;
data_in <= 24'b101100111101001011110011;
#10000;
data_in <= 24'b101101111101011011110111;
#10000;
data_in <= 24'b101111001101100011111010;
#10000;
data_in <= 24'b101011101101000111110011;
#10000;
data_in <= 24'b101011111101000011110001;
#10000;
data_in <= 24'b101011011100111011101111;
#10000;
data_in <= 24'b101100001100111111110000;
#10000;
data_in <= 24'b101101011101010011110101;
#10000;
data_in <= 24'b101110011101100011111001;
#10000;
data_in <= 24'b101110101101100111111010;
#10000;
data_in <= 24'b101110011101100011111001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100011011010001011000001;
#10000;
data_in <= 24'b100101001010110111001101;
#10000;
data_in <= 24'b100111001011011111011001;
#10000;
data_in <= 24'b100111001011100111011110;
#10000;
data_in <= 24'b100101111011011011011101;
#10000;
data_in <= 24'b100100001011001011011101;
#10000;
data_in <= 24'b100010101010110011011010;
#10000;
data_in <= 24'b100001001010100011011000;
#10000;
data_in <= 24'b101000011011100111010111;
#10000;
data_in <= 24'b101010001011111111011111;
#10000;
data_in <= 24'b101010101100001111100101;
#10000;
data_in <= 24'b101001001011111111100100;
#10000;
data_in <= 24'b100111001011100111100000;
#10000;
data_in <= 24'b100100111011001111011110;
#10000;
data_in <= 24'b100011011010111011011100;
#10000;
data_in <= 24'b100010001010100111011010;
#10000;
data_in <= 24'b101101111100111111101101;
#10000;
data_in <= 24'b101110101101000111110001;
#10000;
data_in <= 24'b101101011100111011110000;
#10000;
data_in <= 24'b101010101100010111101010;
#10000;
data_in <= 24'b100111011011101111100100;
#10000;
data_in <= 24'b100101101011010111100010;
#10000;
data_in <= 24'b100100001011000111011111;
#10000;
data_in <= 24'b100011001010110111011110;
#10000;
data_in <= 24'b101111011101011011110110;
#10000;
data_in <= 24'b101111101101011111110111;
#10000;
data_in <= 24'b101110001101001111110101;
#10000;
data_in <= 24'b101011011100100011101101;
#10000;
data_in <= 24'b101000001011111011100111;
#10000;
data_in <= 24'b100101111011100011100101;
#10000;
data_in <= 24'b100100111011010011100010;
#10000;
data_in <= 24'b100011101010111111100000;
#10000;
data_in <= 24'b101111111101100011111000;
#10000;
data_in <= 24'b110000001101100111111001;
#10000;
data_in <= 24'b101110101101010111110111;
#10000;
data_in <= 24'b101011101100101111110000;
#10000;
data_in <= 24'b101000111100000111101010;
#10000;
data_in <= 24'b100110011011101011100111;
#10000;
data_in <= 24'b100100111011010011100010;
#10000;
data_in <= 24'b100011001010110111011110;
#10000;
data_in <= 24'b110000001101110011111011;
#10000;
data_in <= 24'b110000011101110011111110;
#10000;
data_in <= 24'b101111001101100011111011;
#10000;
data_in <= 24'b101100101100111111110100;
#10000;
data_in <= 24'b101001111100010111101110;
#10000;
data_in <= 24'b100111011011110011101001;
#10000;
data_in <= 24'b100100101011001111100001;
#10000;
data_in <= 24'b100010011010101011011100;
#10000;
data_in <= 24'b110000001101110011111011;
#10000;
data_in <= 24'b110000001101101111111101;
#10000;
data_in <= 24'b101111001101100011111011;
#10000;
data_in <= 24'b101100101100111111110110;
#10000;
data_in <= 24'b101010001100011011101111;
#10000;
data_in <= 24'b100111111011111011101011;
#10000;
data_in <= 24'b100101001011010011100101;
#10000;
data_in <= 24'b100010111010101011011101;
#10000;
data_in <= 24'b101111001101100111111000;
#10000;
data_in <= 24'b101111001101100011111010;
#10000;
data_in <= 24'b101101111101010111111000;
#10000;
data_in <= 24'b101011011100110011110011;
#10000;
data_in <= 24'b101001111100010111101110;
#10000;
data_in <= 24'b101000001011111111101100;
#10000;
data_in <= 24'b100101101011011011100111;
#10000;
data_in <= 24'b100011101010110111100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100000001010001111010101;
#10000;
data_in <= 24'b011110001001101111001101;
#10000;
data_in <= 24'b011100011001000111000010;
#10000;
data_in <= 24'b011011011000101110111010;
#10000;
data_in <= 24'b011010111000010110110011;
#10000;
data_in <= 24'b011001000111110110101001;
#10000;
data_in <= 24'b010110000110111010011000;
#10000;
data_in <= 24'b010100010110010010001001;
#10000;
data_in <= 24'b100000011010010011010110;
#10000;
data_in <= 24'b011110011001110011001110;
#10000;
data_in <= 24'b011100111001001011000101;
#10000;
data_in <= 24'b011011101000110010111101;
#10000;
data_in <= 24'b011010101000010110110111;
#10000;
data_in <= 24'b011000110111110110101100;
#10000;
data_in <= 24'b010110000110111110011101;
#10000;
data_in <= 24'b010100010110010010001111;
#10000;
data_in <= 24'b100000101010010111010111;
#10000;
data_in <= 24'b011110111001111011010000;
#10000;
data_in <= 24'b011101011001010011000111;
#10000;
data_in <= 24'b011100001000111010111111;
#10000;
data_in <= 24'b011011001000011110111001;
#10000;
data_in <= 24'b011001010111111110101110;
#10000;
data_in <= 24'b010110110111001010100000;
#10000;
data_in <= 24'b010100110110100110010011;
#10000;
data_in <= 24'b100001001010011111011001;
#10000;
data_in <= 24'b011111111010000011010010;
#10000;
data_in <= 24'b011101111001011011001001;
#10000;
data_in <= 24'b011100101001000011000001;
#10000;
data_in <= 24'b011011101000100110111011;
#10000;
data_in <= 24'b011001111000000110110000;
#10000;
data_in <= 24'b010111010111010110100011;
#10000;
data_in <= 24'b010110000110111010011000;
#10000;
data_in <= 24'b100001111010100011011010;
#10000;
data_in <= 24'b100000011010000111010110;
#10000;
data_in <= 24'b011110011001100011001011;
#10000;
data_in <= 24'b011101001001001011000011;
#10000;
data_in <= 24'b011011111000101010111100;
#10000;
data_in <= 24'b011010001000001010110001;
#10000;
data_in <= 24'b011000000111100010100110;
#10000;
data_in <= 24'b010110100111001010011100;
#10000;
data_in <= 24'b100001111010011111011100;
#10000;
data_in <= 24'b100000101010001011010111;
#10000;
data_in <= 24'b011110111001101011001101;
#10000;
data_in <= 24'b011100111001001011000101;
#10000;
data_in <= 24'b011011101000110010111101;
#10000;
data_in <= 24'b011001111000001110110010;
#10000;
data_in <= 24'b011000000111101010101000;
#10000;
data_in <= 24'b010111000111010110100001;
#10000;
data_in <= 24'b100001111010011111011100;
#10000;
data_in <= 24'b100000101010001011010111;
#10000;
data_in <= 24'b011110111001101011001111;
#10000;
data_in <= 24'b011101001001001111000110;
#10000;
data_in <= 24'b011011101000110010111101;
#10000;
data_in <= 24'b011010001000010010110011;
#10000;
data_in <= 24'b011000000111110110101010;
#10000;
data_in <= 24'b010111000111011110100011;
#10000;
data_in <= 24'b100001111010011111011100;
#10000;
data_in <= 24'b100000101010001011010111;
#10000;
data_in <= 24'b011111001001101111010000;
#10000;
data_in <= 24'b011101001001001111000110;
#10000;
data_in <= 24'b011011101000101110111110;
#10000;
data_in <= 24'b011001101000010010110101;
#10000;
data_in <= 24'b011000000111110010101011;
#10000;
data_in <= 24'b010111010111100010100100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010101010110011110000100;
#10000;
data_in <= 24'b010000000101000101101011;
#10000;
data_in <= 24'b001010100011110101011000;
#10000;
data_in <= 24'b000101110010110001001000;
#10000;
data_in <= 24'b000110000010110101001100;
#10000;
data_in <= 24'b000101110010111101001101;
#10000;
data_in <= 24'b000011110010100101000111;
#10000;
data_in <= 24'b000111110011100101010111;
#10000;
data_in <= 24'b010100110110010010000101;
#10000;
data_in <= 24'b010011000101110001111001;
#10000;
data_in <= 24'b001110010100110101101100;
#10000;
data_in <= 24'b001000000011010101010101;
#10000;
data_in <= 24'b000110100011001101010101;
#10000;
data_in <= 24'b001000010011110101011111;
#10000;
data_in <= 24'b001000100100000101100010;
#10000;
data_in <= 24'b001100110101001001110011;
#10000;
data_in <= 24'b010100010110010010000101;
#10000;
data_in <= 24'b010101000110011010000011;
#10000;
data_in <= 24'b010001110101101101111010;
#10000;
data_in <= 24'b001000100011100101011001;
#10000;
data_in <= 24'b000101100011000101010011;
#10000;
data_in <= 24'b001001010100000101100100;
#10000;
data_in <= 24'b001011110100111101110010;
#10000;
data_in <= 24'b010010000110100010001011;
#10000;
data_in <= 24'b010100010110010110001000;
#10000;
data_in <= 24'b010100110110011110000110;
#10000;
data_in <= 24'b010010100101111101111111;
#10000;
data_in <= 24'b001001110100000001100010;
#10000;
data_in <= 24'b000101100011000001010100;
#10000;
data_in <= 24'b000111000011100101011110;
#10000;
data_in <= 24'b001010010100101101101111;
#10000;
data_in <= 24'b010010100110110010010000;
#10000;
data_in <= 24'b010100010110011110001011;
#10000;
data_in <= 24'b010100000110010010000111;
#10000;
data_in <= 24'b010011100110010010000111;
#10000;
data_in <= 24'b001111000101011001111010;
#10000;
data_in <= 24'b001011110100101001101111;
#10000;
data_in <= 24'b001001000100001101101010;
#10000;
data_in <= 24'b001001110100100001101111;
#10000;
data_in <= 24'b010001010110100110001111;
#10000;
data_in <= 24'b010101000110100110001111;
#10000;
data_in <= 24'b010011100110010010001000;
#10000;
data_in <= 24'b010101010110110110010001;
#10000;
data_in <= 24'b010110010111001110011000;
#10000;
data_in <= 24'b010101110111010010011011;
#10000;
data_in <= 24'b010001010110010110001110;
#10000;
data_in <= 24'b001101010101100010000000;
#10000;
data_in <= 24'b010010000110101110010011;
#10000;
data_in <= 24'b010101110110110110010110;
#10000;
data_in <= 24'b010011010110010010001010;
#10000;
data_in <= 24'b010100100110110010010001;
#10000;
data_in <= 24'b010111010111011110011111;
#10000;
data_in <= 24'b011010101000100010110001;
#10000;
data_in <= 24'b011001011000010110110000;
#10000;
data_in <= 24'b010011010110111110011010;
#10000;
data_in <= 24'b010011110111001010011101;
#10000;
data_in <= 24'b010110010111001010011010;
#10000;
data_in <= 24'b010011000110010110001101;
#10000;
data_in <= 24'b010010000110001010001010;
#10000;
data_in <= 24'b010011100110101010010011;
#10000;
data_in <= 24'b011010001000010110110001;
#10000;
data_in <= 24'b011100011001001110111110;
#10000;
data_in <= 24'b010110110111110010101001;
#10000;
data_in <= 24'b010100110111011010100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000100010010110001000111;
#10000;
data_in <= 24'b001000110011110001010110;
#10000;
data_in <= 24'b001010100100001001011010;
#10000;
data_in <= 24'b001100110100100001011110;
#10000;
data_in <= 24'b001100000100000101010100;
#10000;
data_in <= 24'b001011010011110101001110;
#10000;
data_in <= 24'b010000110101000001100000;
#10000;
data_in <= 24'b010011100101101101101001;
#10000;
data_in <= 24'b010000000101111110000000;
#10000;
data_in <= 24'b001000110100000001011111;
#10000;
data_in <= 24'b000001000001110000111000;
#10000;
data_in <= 24'b000011000010001000111011;
#10000;
data_in <= 24'b001000000011000101000110;
#10000;
data_in <= 24'b001010110011100101001011;
#10000;
data_in <= 24'b010011010101011101101000;
#10000;
data_in <= 24'b011000110110111001111100;
#10000;
data_in <= 24'b011101001001010010110111;
#10000;
data_in <= 24'b010010010110100010001001;
#10000;
data_in <= 24'b000011000010011001000100;
#10000;
data_in <= 24'b000000110001101000110100;
#10000;
data_in <= 24'b000111110011010001001010;
#10000;
data_in <= 24'b001111000100110101100000;
#10000;
data_in <= 24'b010110110110100101111011;
#10000;
data_in <= 24'b011001110111010010000100;
#10000;
data_in <= 24'b100010011010101111001111;
#10000;
data_in <= 24'b100000111010001111000110;
#10000;
data_in <= 24'b010000110110000001111111;
#10000;
data_in <= 24'b000011000010011001000100;
#10000;
data_in <= 24'b000101100010101101000110;
#10000;
data_in <= 24'b001110110101000001100110;
#10000;
data_in <= 24'b010101110110100001111101;
#10000;
data_in <= 24'b010100100110000101110100;
#10000;
data_in <= 24'b100001101010101011010000;
#10000;
data_in <= 24'b101001001100011011101010;
#10000;
data_in <= 24'b011011111000110110110000;
#10000;
data_in <= 24'b000110010011010101010100;
#10000;
data_in <= 24'b000000000001010000110010;
#10000;
data_in <= 24'b000011110010011001000000;
#10000;
data_in <= 24'b001011000100000001011001;
#10000;
data_in <= 24'b001100000100010001011101;
#10000;
data_in <= 24'b011110101001110111000101;
#10000;
data_in <= 24'b101000011100010111101011;
#10000;
data_in <= 24'b100001011010010111001001;
#10000;
data_in <= 24'b010000100110000010000011;
#10000;
data_in <= 24'b000100010010110001001110;
#10000;
data_in <= 24'b000000000000111000101100;
#10000;
data_in <= 24'b000000000001010000110011;
#10000;
data_in <= 24'b000101000010101001000110;
#10000;
data_in <= 24'b011100001001001110111110;
#10000;
data_in <= 24'b100101001011011111011111;
#10000;
data_in <= 24'b100010111010101111010100;
#10000;
data_in <= 24'b011100101001000110111000;
#10000;
data_in <= 24'b010011110110101010001111;
#10000;
data_in <= 24'b000011110010101001001100;
#10000;
data_in <= 24'b000000000000110000101110;
#10000;
data_in <= 24'b000000010001100000111000;
#10000;
data_in <= 24'b011011111001001010111101;
#10000;
data_in <= 24'b100011001010111011011001;
#10000;
data_in <= 24'b100001001010010011001101;
#10000;
data_in <= 24'b100000001001111111000110;
#10000;
data_in <= 24'b011100101000111110110100;
#10000;
data_in <= 24'b001100010100110001110001;
#10000;
data_in <= 24'b000000000001100000111100;
#10000;
data_in <= 24'b000000000001001000110100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001110100100110101100010;
#10000;
data_in <= 24'b001100010100011001011100;
#10000;
data_in <= 24'b001100000100010001011101;
#10000;
data_in <= 24'b000110100011000001001100;
#10000;
data_in <= 24'b000110100011001001010000;
#10000;
data_in <= 24'b001111010101100001111010;
#10000;
data_in <= 24'b010101110111001110010110;
#10000;
data_in <= 24'b011001000111111110100100;
#10000;
data_in <= 24'b001011000011111101010100;
#10000;
data_in <= 24'b001010110011110101010100;
#10000;
data_in <= 24'b001100010100010101011110;
#10000;
data_in <= 24'b000111100011010001010000;
#10000;
data_in <= 24'b000110110011001101010001;
#10000;
data_in <= 24'b001110110101010001110110;
#10000;
data_in <= 24'b010101000110111010010010;
#10000;
data_in <= 24'b011000100111110110100010;
#10000;
data_in <= 24'b000111110011000001000101;
#10000;
data_in <= 24'b001000110011010101001100;
#10000;
data_in <= 24'b001100000100010001011101;
#10000;
data_in <= 24'b001001000011100101010100;
#10000;
data_in <= 24'b000111100011001101010010;
#10000;
data_in <= 24'b001101100100111101110001;
#10000;
data_in <= 24'b010011100110100010001100;
#10000;
data_in <= 24'b011000000111110010011111;
#10000;
data_in <= 24'b000111000010110101000010;
#10000;
data_in <= 24'b000111110011001001000111;
#10000;
data_in <= 24'b001100000100000101011011;
#10000;
data_in <= 24'b001001000011100101010100;
#10000;
data_in <= 24'b000111010011001001010001;
#10000;
data_in <= 24'b001100010100101001101010;
#10000;
data_in <= 24'b010010000110001110000101;
#10000;
data_in <= 24'b010111010111100110011100;
#10000;
data_in <= 24'b001000010011001001000111;
#10000;
data_in <= 24'b000111100011000101000110;
#10000;
data_in <= 24'b001011000011110101010111;
#10000;
data_in <= 24'b001000010011011001010001;
#10000;
data_in <= 24'b000110010010111101001011;
#10000;
data_in <= 24'b001010100100001101100011;
#10000;
data_in <= 24'b010000010101110001111110;
#10000;
data_in <= 24'b010110000111001010010110;
#10000;
data_in <= 24'b001000000011000101000110;
#10000;
data_in <= 24'b000111000010111101000100;
#10000;
data_in <= 24'b001010100011110001010011;
#10000;
data_in <= 24'b001000000011010101010000;
#10000;
data_in <= 24'b000101010010101101000111;
#10000;
data_in <= 24'b001000000011100101011001;
#10000;
data_in <= 24'b001101110101000001110010;
#10000;
data_in <= 24'b010011110110100110001101;
#10000;
data_in <= 24'b000101000010010100111000;
#10000;
data_in <= 24'b000101010010100000111101;
#10000;
data_in <= 24'b001010100011110001010011;
#10000;
data_in <= 24'b001000100011011101010010;
#10000;
data_in <= 24'b000100010010011101000011;
#10000;
data_in <= 24'b000101010010111001001110;
#10000;
data_in <= 24'b001010100100001101100101;
#10000;
data_in <= 24'b010000110101110110000001;
#10000;
data_in <= 24'b000010010001100100101010;
#10000;
data_in <= 24'b000100000010000100110100;
#10000;
data_in <= 24'b001010110011111001010011;
#10000;
data_in <= 24'b001001110011110001010010;
#10000;
data_in <= 24'b000100010010011001000001;
#10000;
data_in <= 24'b000100000010011001000010;
#10000;
data_in <= 24'b001000100011100101011001;
#10000;
data_in <= 24'b001111010101011001111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000100111111110100110;
#10000;
data_in <= 24'b010111100111101110100010;
#10000;
data_in <= 24'b010100010110110010010001;
#10000;
data_in <= 24'b010000010101101101111111;
#10000;
data_in <= 24'b010000010101100101111101;
#10000;
data_in <= 24'b010001110101110110000000;
#10000;
data_in <= 24'b001111010101001001110010;
#10000;
data_in <= 24'b001010100011111001011101;
#10000;
data_in <= 24'b011000111000000010100111;
#10000;
data_in <= 24'b010110100111010110011010;
#10000;
data_in <= 24'b010011010110011110001100;
#10000;
data_in <= 24'b010001000101110010000000;
#10000;
data_in <= 24'b001111110101010101111000;
#10000;
data_in <= 24'b001111000101000101110001;
#10000;
data_in <= 24'b001101110100101101101010;
#10000;
data_in <= 24'b001101010100011101100110;
#10000;
data_in <= 24'b011001111000001010100111;
#10000;
data_in <= 24'b010110000111001110011000;
#10000;
data_in <= 24'b010010110110010110001010;
#10000;
data_in <= 24'b010001010101110110000001;
#10000;
data_in <= 24'b001110100101000001110011;
#10000;
data_in <= 24'b001100000100010101100101;
#10000;
data_in <= 24'b001101010100100101101000;
#10000;
data_in <= 24'b010001000101011001110101;
#10000;
data_in <= 24'b011001011000000010100101;
#10000;
data_in <= 24'b010111000111011110011100;
#10000;
data_in <= 24'b010100010110101110001111;
#10000;
data_in <= 24'b010001010101111010000000;
#10000;
data_in <= 24'b001101110100110101110000;
#10000;
data_in <= 24'b001100010100011001100110;
#10000;
data_in <= 24'b001111100101001001110001;
#10000;
data_in <= 24'b010100100110010010000011;
#10000;
data_in <= 24'b010111100111100110011110;
#10000;
data_in <= 24'b011000000111101110100000;
#10000;
data_in <= 24'b010101110111000110010101;
#10000;
data_in <= 24'b010000010101101001111100;
#10000;
data_in <= 24'b001100110100100101101100;
#10000;
data_in <= 24'b001110100100111101101111;
#10000;
data_in <= 24'b010010100101111001111101;
#10000;
data_in <= 24'b010101100110100010000111;
#10000;
data_in <= 24'b010101110111001010010111;
#10000;
data_in <= 24'b011000000111101110100000;
#10000;
data_in <= 24'b010101100111000010010100;
#10000;
data_in <= 24'b001110110101010001110110;
#10000;
data_in <= 24'b001100100100100001101011;
#10000;
data_in <= 24'b010000110101100001111000;
#10000;
data_in <= 24'b010100010110001110000010;
#10000;
data_in <= 24'b010100010110000101111110;
#10000;
data_in <= 24'b010101010111000010010101;
#10000;
data_in <= 24'b010111000111011110011100;
#10000;
data_in <= 24'b010100000110101010001110;
#10000;
data_in <= 24'b001110010101001001110100;
#10000;
data_in <= 24'b001101100100110001101111;
#10000;
data_in <= 24'b010001110101110001111100;
#10000;
data_in <= 24'b010011110110000110000000;
#10000;
data_in <= 24'b010001100101011001110011;
#10000;
data_in <= 24'b010110110111010010010110;
#10000;
data_in <= 24'b010110110111001110010111;
#10000;
data_in <= 24'b010011100110011110001001;
#10000;
data_in <= 24'b001111010101001101110110;
#10000;
data_in <= 24'b001111010101001001110010;
#10000;
data_in <= 24'b010010010101111001111110;
#10000;
data_in <= 24'b010010010101110101111100;
#10000;
data_in <= 24'b010000000101000001101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001001010011011101010110;
#10000;
data_in <= 24'b001111010100110001101100;
#10000;
data_in <= 24'b010011010101101001111010;
#10000;
data_in <= 24'b010010000101011001110011;
#10000;
data_in <= 24'b001111100100110001101001;
#10000;
data_in <= 24'b001110110100100101100101;
#10000;
data_in <= 24'b001111100100100101100111;
#10000;
data_in <= 24'b001110110100100101100110;
#10000;
data_in <= 24'b010010000101011101110111;
#10000;
data_in <= 24'b010011100101111001111011;
#10000;
data_in <= 24'b010100000101111001111011;
#10000;
data_in <= 24'b010001010101001101101111;
#10000;
data_in <= 24'b001110100100011001100010;
#10000;
data_in <= 24'b001101100100001101011101;
#10000;
data_in <= 24'b001101110100010001011110;
#10000;
data_in <= 24'b001110000100010101011111;
#10000;
data_in <= 24'b010101010110010110000010;
#10000;
data_in <= 24'b010100000101111001111011;
#10000;
data_in <= 24'b010010010101010001110010;
#10000;
data_in <= 24'b010000000100110001101000;
#10000;
data_in <= 24'b001101110100001001011101;
#10000;
data_in <= 24'b001100100011111001010110;
#10000;
data_in <= 24'b001101010100001001011000;
#10000;
data_in <= 24'b001111010100101001100000;
#10000;
data_in <= 24'b010011100101110001111001;
#10000;
data_in <= 24'b010000110101000101101101;
#10000;
data_in <= 24'b001111000100100001100100;
#10000;
data_in <= 24'b001110010100011001100000;
#10000;
data_in <= 24'b001101000100000001011000;
#10000;
data_in <= 24'b001011010011101001010000;
#10000;
data_in <= 24'b001101100100000101010101;
#10000;
data_in <= 24'b010001000101000001100010;
#10000;
data_in <= 24'b010011000101101001110111;
#10000;
data_in <= 24'b010000010100110101101001;
#10000;
data_in <= 24'b001110000100001101011110;
#10000;
data_in <= 24'b001101000100000001011000;
#10000;
data_in <= 24'b001011110011101001001110;
#10000;
data_in <= 24'b001010100011011001001000;
#10000;
data_in <= 24'b001110000100001001010011;
#10000;
data_in <= 24'b010010110101010101100110;
#10000;
data_in <= 24'b010010100101100001110100;
#10000;
data_in <= 24'b001111110100110001100110;
#10000;
data_in <= 24'b001100110011111101010111;
#10000;
data_in <= 24'b001011010011101001010000;
#10000;
data_in <= 24'b001010100011011001001000;
#10000;
data_in <= 24'b001011000011100101001001;
#10000;
data_in <= 24'b010000000100101101011001;
#10000;
data_in <= 24'b010101010110000101101101;
#10000;
data_in <= 24'b010000110101000001101010;
#10000;
data_in <= 24'b001110000100010001011100;
#10000;
data_in <= 24'b001011100011100101001111;
#10000;
data_in <= 24'b001010010011010001001000;
#10000;
data_in <= 24'b001011000011011001000111;
#10000;
data_in <= 24'b001101000011111101001101;
#10000;
data_in <= 24'b010001010100111001011011;
#10000;
data_in <= 24'b010101000101111001101000;
#10000;
data_in <= 24'b001111010100101101100010;
#10000;
data_in <= 24'b001101100100000101010111;
#10000;
data_in <= 24'b001010110011011001001010;
#10000;
data_in <= 24'b001010010011001101000100;
#10000;
data_in <= 24'b001011010011100001000110;
#10000;
data_in <= 24'b001101100100000001001010;
#10000;
data_in <= 24'b001111010100011001010000;
#10000;
data_in <= 24'b010000000100101101010011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001110100100100001100101;
#10000;
data_in <= 24'b010000010101000001110000;
#10000;
data_in <= 24'b010000100101001101110100;
#10000;
data_in <= 24'b010001110101101001111101;
#10000;
data_in <= 24'b010101000110011010001011;
#10000;
data_in <= 24'b010110100110110110010011;
#10000;
data_in <= 24'b010111110111010010011010;
#10000;
data_in <= 24'b011010011000000010100110;
#10000;
data_in <= 24'b010001000101000001101100;
#10000;
data_in <= 24'b010011010101101101110111;
#10000;
data_in <= 24'b010100000101111101111111;
#10000;
data_in <= 24'b010100110110010010000101;
#10000;
data_in <= 24'b010110110110101110001111;
#10000;
data_in <= 24'b010110110110110110010010;
#10000;
data_in <= 24'b010111010111000010010101;
#10000;
data_in <= 24'b011001110111101010011111;
#10000;
data_in <= 24'b010010110101011101101111;
#10000;
data_in <= 24'b010101100110010001111011;
#10000;
data_in <= 24'b010110110110011110000011;
#10000;
data_in <= 24'b010110100110100010000101;
#10000;
data_in <= 24'b010111010110110010001100;
#10000;
data_in <= 24'b010111100110111110010000;
#10000;
data_in <= 24'b011001000111010010011000;
#10000;
data_in <= 24'b011011101000000110100100;
#10000;
data_in <= 24'b010110010110010001111000;
#10000;
data_in <= 24'b011010000111010110001011;
#10000;
data_in <= 24'b011100010111110110010101;
#10000;
data_in <= 24'b011100000111110110010111;
#10000;
data_in <= 24'b011011110111110110011010;
#10000;
data_in <= 24'b011010010111100010011000;
#10000;
data_in <= 24'b011010000111011110011000;
#10000;
data_in <= 24'b011011010111111010011111;
#10000;
data_in <= 24'b011001010110111110000000;
#10000;
data_in <= 24'b011101011000000110010011;
#10000;
data_in <= 24'b011110101000100010011011;
#10000;
data_in <= 24'b011100000111111010010100;
#10000;
data_in <= 24'b011001000111000110001011;
#10000;
data_in <= 24'b010011110101110101111001;
#10000;
data_in <= 24'b001111110100110101101010;
#10000;
data_in <= 24'b001110010100100001101000;
#10000;
data_in <= 24'b011101011000000010001110;
#10000;
data_in <= 24'b011101111000001010010000;
#10000;
data_in <= 24'b011000100110111010000000;
#10000;
data_in <= 24'b010000010100111101100010;
#10000;
data_in <= 24'b001011100011101001010010;
#10000;
data_in <= 24'b001000010010111001001000;
#10000;
data_in <= 24'b000111000010100001000100;
#10000;
data_in <= 24'b000110110010101001001010;
#10000;
data_in <= 24'b011010000111010010000000;
#10000;
data_in <= 24'b010111000110100001110100;
#10000;
data_in <= 24'b001101100100001101010011;
#10000;
data_in <= 24'b000011110001110100101111;
#10000;
data_in <= 24'b000010110001100000101110;
#10000;
data_in <= 24'b000111010010101101000010;
#10000;
data_in <= 24'b001110010100010101100001;
#10000;
data_in <= 24'b010011010101101101111000;
#10000;
data_in <= 24'b001011010011011101000001;
#10000;
data_in <= 24'b001000110010111100111011;
#10000;
data_in <= 24'b000001010001001000100000;
#10000;
data_in <= 24'b000000000000000000001110;
#10000;
data_in <= 24'b000000010000111000100100;
#10000;
data_in <= 24'b001011000011100101010011;
#10000;
data_in <= 24'b010110000110011010000011;
#10000;
data_in <= 24'b011101101000010110100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011100111000100110101101;
#10000;
data_in <= 24'b011100011000100110101101;
#10000;
data_in <= 24'b011100111000110110110001;
#10000;
data_in <= 24'b011111011001100110111100;
#10000;
data_in <= 24'b100001101010011011001010;
#10000;
data_in <= 24'b100100001011001011010110;
#10000;
data_in <= 24'b100101111011110111100000;
#10000;
data_in <= 24'b100110101100001011100101;
#10000;
data_in <= 24'b011011111000010110101001;
#10000;
data_in <= 24'b011111011001010110111001;
#10000;
data_in <= 24'b100011001010010011001000;
#10000;
data_in <= 24'b100011101010101011001101;
#10000;
data_in <= 24'b100010011010100111001101;
#10000;
data_in <= 24'b100010011010110111010001;
#10000;
data_in <= 24'b100100011011011111011010;
#10000;
data_in <= 24'b100100111011110111100010;
#10000;
data_in <= 24'b100001001001100010111011;
#10000;
data_in <= 24'b100110001011000111010011;
#10000;
data_in <= 24'b101001101011111011100010;
#10000;
data_in <= 24'b100110101011011011011001;
#10000;
data_in <= 24'b100011001010110011010000;
#10000;
data_in <= 24'b100010111010111111010101;
#10000;
data_in <= 24'b100101001011100111011111;
#10000;
data_in <= 24'b100101001011110111100100;
#10000;
data_in <= 24'b011101001000100010101011;
#10000;
data_in <= 24'b100100101010100011001011;
#10000;
data_in <= 24'b101001011011110111100001;
#10000;
data_in <= 24'b100111011011100111011100;
#10000;
data_in <= 24'b100100101011000111011000;
#10000;
data_in <= 24'b100101001011100011011110;
#10000;
data_in <= 24'b100101101011101011100010;
#10000;
data_in <= 24'b100100001011011111011110;
#10000;
data_in <= 24'b001101110100101001101011;
#10000;
data_in <= 24'b011010010111111110100010;
#10000;
data_in <= 24'b100101111010111111010011;
#10000;
data_in <= 24'b100111111011101111011110;
#10000;
data_in <= 24'b100101111011011011011101;
#10000;
data_in <= 24'b100101011011100111011111;
#10000;
data_in <= 24'b100100011011010111011101;
#10000;
data_in <= 24'b100001101010110011010110;
#10000;
data_in <= 24'b001100100100010101100110;
#10000;
data_in <= 24'b011010010111111110100010;
#10000;
data_in <= 24'b100110111011001111010111;
#10000;
data_in <= 24'b101000101011111011100001;
#10000;
data_in <= 24'b100100111011001011011001;
#10000;
data_in <= 24'b100011011011000111010111;
#10000;
data_in <= 24'b100100001011001111011110;
#10000;
data_in <= 24'b100011101011010011011110;
#10000;
data_in <= 24'b011010100111110110011110;
#10000;
data_in <= 24'b100010101010000011000011;
#10000;
data_in <= 24'b101001101011111011100010;
#10000;
data_in <= 24'b101000111011111111100010;
#10000;
data_in <= 24'b100101001011001111011010;
#10000;
data_in <= 24'b100011101011001011011000;
#10000;
data_in <= 24'b100100011011010011011111;
#10000;
data_in <= 24'b100100001011011011100000;
#10000;
data_in <= 24'b100010101001111110111110;
#10000;
data_in <= 24'b100110001010111111001111;
#10000;
data_in <= 24'b101000011011110011011110;
#10000;
data_in <= 24'b101000011011111111100010;
#10000;
data_in <= 24'b100111101011111011100010;
#10000;
data_in <= 24'b100110001011110011100010;
#10000;
data_in <= 24'b100010111011001011011001;
#10000;
data_in <= 24'b011111011010010111001111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101000101100110011110001;
#10000;
data_in <= 24'b101000001100110011110001;
#10000;
data_in <= 24'b101000001100110011110001;
#10000;
data_in <= 24'b100111011100100111101110;
#10000;
data_in <= 24'b100101011100000111100110;
#10000;
data_in <= 24'b100010111011011111011100;
#10000;
data_in <= 24'b100001101011001011010111;
#10000;
data_in <= 24'b100001001011000011010101;
#10000;
data_in <= 24'b100111011100011111101100;
#10000;
data_in <= 24'b100111011100100111101110;
#10000;
data_in <= 24'b100111111100101111110000;
#10000;
data_in <= 24'b100111001100100011101101;
#10000;
data_in <= 24'b100101011100000111100110;
#10000;
data_in <= 24'b100011001011100011011101;
#10000;
data_in <= 24'b100001101011001011010111;
#10000;
data_in <= 24'b100000111010111011010101;
#10000;
data_in <= 24'b100110011100001011101001;
#10000;
data_in <= 24'b100110111100011011101101;
#10000;
data_in <= 24'b100111111100101011110001;
#10000;
data_in <= 24'b100111101100100111110000;
#10000;
data_in <= 24'b100110111100010111101010;
#10000;
data_in <= 24'b100100111011110111100010;
#10000;
data_in <= 24'b100010111011010111011010;
#10000;
data_in <= 24'b100001101010111111010110;
#10000;
data_in <= 24'b100101011011111011100101;
#10000;
data_in <= 24'b100110011100010011101011;
#10000;
data_in <= 24'b100111111100101011110001;
#10000;
data_in <= 24'b101000101100101111110010;
#10000;
data_in <= 24'b101000001100101011101111;
#10000;
data_in <= 24'b100111011100010011101010;
#10000;
data_in <= 24'b100101111011110011100010;
#10000;
data_in <= 24'b100011101011010111011100;
#10000;
data_in <= 24'b100100001011100011100010;
#10000;
data_in <= 24'b100110001100000011101010;
#10000;
data_in <= 24'b100111111100011111110001;
#10000;
data_in <= 24'b101000111100101011110001;
#10000;
data_in <= 24'b101001101100101111110001;
#10000;
data_in <= 24'b101001011100101011110000;
#10000;
data_in <= 24'b100111111100001111100111;
#10000;
data_in <= 24'b100101111011101111100001;
#10000;
data_in <= 24'b100010111011001111011101;
#10000;
data_in <= 24'b100100111011101111100101;
#10000;
data_in <= 24'b100111001100001011101100;
#10000;
data_in <= 24'b101000011100010111101101;
#10000;
data_in <= 24'b101001101100100111110001;
#10000;
data_in <= 24'b101011001100110111110100;
#10000;
data_in <= 24'b101010001100101011101110;
#10000;
data_in <= 24'b100111111100000011100111;
#10000;
data_in <= 24'b100010001010111111011011;
#10000;
data_in <= 24'b100100011011100011100100;
#10000;
data_in <= 24'b100110011011111111101001;
#10000;
data_in <= 24'b100111101100001011101010;
#10000;
data_in <= 24'b101001101100100111110001;
#10000;
data_in <= 24'b101100001101000111111000;
#10000;
data_in <= 24'b101100011101000111110101;
#10000;
data_in <= 24'b101010011100100011101111;
#10000;
data_in <= 24'b100010011011000011011100;
#10000;
data_in <= 24'b100100011011100011100100;
#10000;
data_in <= 24'b100110011011111111101001;
#10000;
data_in <= 24'b100111101100001011101010;
#10000;
data_in <= 24'b101001111100101111110001;
#10000;
data_in <= 24'b101101001101011011111010;
#10000;
data_in <= 24'b101110001101010111111010;
#10000;
data_in <= 24'b101100011100111011110101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100010001011001111011010;
#10000;
data_in <= 24'b100010111011011011011101;
#10000;
data_in <= 24'b100100001011101011100100;
#10000;
data_in <= 24'b100101111100000011100111;
#10000;
data_in <= 24'b100110111100010011101011;
#10000;
data_in <= 24'b100111011100011011101101;
#10000;
data_in <= 24'b101000001100011111101110;
#10000;
data_in <= 24'b101000101100011111101101;
#10000;
data_in <= 24'b100001101011000011011010;
#10000;
data_in <= 24'b100010001011001011011100;
#10000;
data_in <= 24'b100011001011011011100000;
#10000;
data_in <= 24'b100100011011101111100101;
#10000;
data_in <= 24'b100101011011111111101001;
#10000;
data_in <= 24'b100110111100001111101101;
#10000;
data_in <= 24'b100111101100011011110000;
#10000;
data_in <= 24'b101000011100100011101111;
#10000;
data_in <= 24'b100001011010110111010111;
#10000;
data_in <= 24'b100001101010110111011001;
#10000;
data_in <= 24'b100010001010111111011011;
#10000;
data_in <= 24'b100010111011001011011110;
#10000;
data_in <= 24'b100100001011011111100011;
#10000;
data_in <= 24'b100101101011111011101000;
#10000;
data_in <= 24'b100110111100001111101101;
#10000;
data_in <= 24'b100111101100011111101110;
#10000;
data_in <= 24'b100001111010110111010111;
#10000;
data_in <= 24'b100001011010101011010110;
#10000;
data_in <= 24'b100001011010101011010110;
#10000;
data_in <= 24'b100001001010101111010111;
#10000;
data_in <= 24'b100010011011000011011100;
#10000;
data_in <= 24'b100100001011011111100011;
#10000;
data_in <= 24'b100101111011111011101010;
#10000;
data_in <= 24'b100111001100010011101110;
#10000;
data_in <= 24'b100100001011001011011101;
#10000;
data_in <= 24'b100011001010111111011011;
#10000;
data_in <= 24'b100010001010101011011000;
#10000;
data_in <= 24'b100001001010100011010110;
#10000;
data_in <= 24'b100001111010101111011001;
#10000;
data_in <= 24'b100011011011001011011110;
#10000;
data_in <= 24'b100101011011101011100110;
#10000;
data_in <= 24'b100110101100000011101010;
#10000;
data_in <= 24'b100110111011101111100110;
#10000;
data_in <= 24'b100101001011010111100010;
#10000;
data_in <= 24'b100011011010111011011100;
#10000;
data_in <= 24'b100001111010100111010111;
#10000;
data_in <= 24'b100001111010100111010111;
#10000;
data_in <= 24'b100010011010110111011011;
#10000;
data_in <= 24'b100011111011010011100000;
#10000;
data_in <= 24'b100101001011101011100100;
#10000;
data_in <= 24'b101000111100000011101100;
#10000;
data_in <= 24'b100111001011100111100110;
#10000;
data_in <= 24'b100100101010111011011101;
#10000;
data_in <= 24'b100010001010011011010101;
#10000;
data_in <= 24'b100000101010001111010001;
#10000;
data_in <= 24'b100000111010010111010011;
#10000;
data_in <= 24'b100010001010101111010111;
#10000;
data_in <= 24'b100010111010111011011001;
#10000;
data_in <= 24'b101001011100000011101100;
#10000;
data_in <= 24'b100111001011100111100110;
#10000;
data_in <= 24'b100100011010110111011100;
#10000;
data_in <= 24'b100001001010001011010001;
#10000;
data_in <= 24'b011111111001110111001100;
#10000;
data_in <= 24'b011111011001111011001100;
#10000;
data_in <= 24'b100000001010000111001110;
#10000;
data_in <= 24'b100000111010010011010001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101001101100101011101110;
#10000;
data_in <= 24'b101001111100110011101110;
#10000;
data_in <= 24'b101011001100111111110001;
#10000;
data_in <= 24'b101100111101001111110110;
#10000;
data_in <= 24'b101101111101100011111001;
#10000;
data_in <= 24'b101110001101100111111010;
#10000;
data_in <= 24'b101110011101100011110111;
#10000;
data_in <= 24'b101110011101100011110111;
#10000;
data_in <= 24'b101001011100101011110000;
#10000;
data_in <= 24'b101001101100110011101111;
#10000;
data_in <= 24'b101010111101000011110010;
#10000;
data_in <= 24'b101100011101010011110110;
#10000;
data_in <= 24'b101101111101100011111001;
#10000;
data_in <= 24'b101110001101101011111000;
#10000;
data_in <= 24'b101110101101100111111000;
#10000;
data_in <= 24'b101110011101100011110111;
#10000;
data_in <= 24'b101000111100101011110000;
#10000;
data_in <= 24'b101001111100110111110000;
#10000;
data_in <= 24'b101010111101000011110010;
#10000;
data_in <= 24'b101100001101001111110101;
#10000;
data_in <= 24'b101101001101010111110110;
#10000;
data_in <= 24'b101101101101100011110110;
#10000;
data_in <= 24'b101110001101100011110101;
#10000;
data_in <= 24'b101101111101011111110100;
#10000;
data_in <= 24'b101000101100100111110000;
#10000;
data_in <= 24'b101010011100111111110010;
#10000;
data_in <= 24'b101011011101001011110100;
#10000;
data_in <= 24'b101011111101001011110011;
#10000;
data_in <= 24'b101100101101010011110010;
#10000;
data_in <= 24'b101101001101011011110011;
#10000;
data_in <= 24'b101101101101011111110001;
#10000;
data_in <= 24'b101101001101010111101111;
#10000;
data_in <= 24'b101001001100100011110000;
#10000;
data_in <= 24'b101010111101000111110100;
#10000;
data_in <= 24'b101100011101011011111000;
#10000;
data_in <= 24'b101100101101010111110110;
#10000;
data_in <= 24'b101100111101010111110010;
#10000;
data_in <= 24'b101101101101011111110001;
#10000;
data_in <= 24'b101101111101011011101111;
#10000;
data_in <= 24'b101100101101001111101101;
#10000;
data_in <= 24'b101000001100010011101100;
#10000;
data_in <= 24'b101010101101000011110011;
#10000;
data_in <= 24'b101101001101011111111001;
#10000;
data_in <= 24'b101100111101011111110101;
#10000;
data_in <= 24'b101101101101011011110011;
#10000;
data_in <= 24'b101110001101101011110010;
#10000;
data_in <= 24'b101110011101100111110000;
#10000;
data_in <= 24'b101100101101010011101100;
#10000;
data_in <= 24'b100101001011100011100000;
#10000;
data_in <= 24'b101000101100100011101011;
#10000;
data_in <= 24'b101011111101001011110100;
#10000;
data_in <= 24'b101011111101001111110001;
#10000;
data_in <= 24'b101101001101010111101111;
#10000;
data_in <= 24'b101101111101100111110001;
#10000;
data_in <= 24'b101110001101100011101111;
#10000;
data_in <= 24'b101100111101001011101011;
#10000;
data_in <= 24'b100010101010110111010101;
#10000;
data_in <= 24'b100110101011111011100100;
#10000;
data_in <= 24'b101010001100101011101110;
#10000;
data_in <= 24'b101011001100110111101110;
#10000;
data_in <= 24'b101100001101000011101101;
#10000;
data_in <= 24'b101101001101010111101111;
#10000;
data_in <= 24'b101101011101010011101101;
#10000;
data_in <= 24'b101100001100111011101001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101111001101101111111100;
#10000;
data_in <= 24'b101110011101100011111001;
#10000;
data_in <= 24'b101100111101000111110100;
#10000;
data_in <= 24'b101010111100101011110001;
#10000;
data_in <= 24'b101001101100001111101111;
#10000;
data_in <= 24'b100111111011110111101100;
#10000;
data_in <= 24'b100101111011011111101000;
#10000;
data_in <= 24'b100100111011001011100101;
#10000;
data_in <= 24'b101110011101100011111001;
#10000;
data_in <= 24'b101101101101010011110111;
#10000;
data_in <= 24'b101100011100111011110011;
#10000;
data_in <= 24'b101010011100100011101111;
#10000;
data_in <= 24'b101000101100001011101101;
#10000;
data_in <= 24'b100111001011101011101001;
#10000;
data_in <= 24'b100101011011010111100110;
#10000;
data_in <= 24'b100100011011000011100101;
#10000;
data_in <= 24'b101101001101011011110100;
#10000;
data_in <= 24'b101100001101000011110011;
#10000;
data_in <= 24'b101010111100101111101111;
#10000;
data_in <= 24'b101001101100010011101101;
#10000;
data_in <= 24'b100111111011111111101010;
#10000;
data_in <= 24'b100110011011011111100110;
#10000;
data_in <= 24'b100100101011000111100100;
#10000;
data_in <= 24'b100011101010110111100010;
#10000;
data_in <= 24'b101100011101001111110001;
#10000;
data_in <= 24'b101011101100111011110001;
#10000;
data_in <= 24'b101010011100100111101101;
#10000;
data_in <= 24'b101001011100001111101100;
#10000;
data_in <= 24'b100111101011111011101001;
#10000;
data_in <= 24'b100110001011011011100101;
#10000;
data_in <= 24'b100100001010111111100010;
#10000;
data_in <= 24'b100011001010101111100000;
#10000;
data_in <= 24'b101011111101000111101111;
#10000;
data_in <= 24'b101010101100110111101111;
#10000;
data_in <= 24'b101001101100100011101100;
#10000;
data_in <= 24'b101000101100001011101011;
#10000;
data_in <= 24'b100111101011110111101010;
#10000;
data_in <= 24'b100110001011011011100111;
#10000;
data_in <= 24'b100100011010111011100001;
#10000;
data_in <= 24'b100011011010100111011111;
#10000;
data_in <= 24'b101011011100111111101101;
#10000;
data_in <= 24'b101010011100110011101110;
#10000;
data_in <= 24'b101001101100100011101100;
#10000;
data_in <= 24'b101000101100001011101011;
#10000;
data_in <= 24'b100111011011110011101001;
#10000;
data_in <= 24'b100101111011010111100110;
#10000;
data_in <= 24'b100100001010110111100000;
#10000;
data_in <= 24'b100011001010100011011110;
#10000;
data_in <= 24'b101010111100110111101011;
#10000;
data_in <= 24'b101001111100101011101100;
#10000;
data_in <= 24'b101001001100011011101010;
#10000;
data_in <= 24'b101000011100000111101010;
#10000;
data_in <= 24'b100111001011101111101000;
#10000;
data_in <= 24'b100101101011010011100101;
#10000;
data_in <= 24'b100011111010110011011111;
#10000;
data_in <= 24'b100010101010011011011100;
#10000;
data_in <= 24'b101010011100101011101011;
#10000;
data_in <= 24'b101001011100011111101011;
#10000;
data_in <= 24'b101000111100010011101011;
#10000;
data_in <= 24'b101000001100000011101001;
#10000;
data_in <= 24'b100110111011101011100111;
#10000;
data_in <= 24'b100101011011001111100100;
#10000;
data_in <= 24'b100011101010101111011110;
#10000;
data_in <= 24'b100001111010011011011011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100010111010101011011111;
#10000;
data_in <= 24'b100001011010001111011010;
#10000;
data_in <= 24'b011111001001101111010000;
#10000;
data_in <= 24'b011100101001000111000100;
#10000;
data_in <= 24'b011010111000101010111101;
#10000;
data_in <= 24'b011001001000010010110101;
#10000;
data_in <= 24'b011000010111111110101110;
#10000;
data_in <= 24'b011000000111110110101010;
#10000;
data_in <= 24'b100010111010100111100000;
#10000;
data_in <= 24'b100001011010001111011010;
#10000;
data_in <= 24'b011110111001101011001111;
#10000;
data_in <= 24'b011100101001000111000110;
#10000;
data_in <= 24'b011010101000100110111100;
#10000;
data_in <= 24'b011000111000001110110100;
#10000;
data_in <= 24'b011000000111111010101101;
#10000;
data_in <= 24'b010111110111110010101001;
#10000;
data_in <= 24'b100010011010011111011110;
#10000;
data_in <= 24'b100000111010000111011000;
#10000;
data_in <= 24'b011110101001100111001110;
#10000;
data_in <= 24'b011100011001000011000101;
#10000;
data_in <= 24'b011010011000100010111011;
#10000;
data_in <= 24'b011000101000001010110011;
#10000;
data_in <= 24'b010111010111111010101100;
#10000;
data_in <= 24'b010111000111101010101001;
#10000;
data_in <= 24'b100010001010011011011101;
#10000;
data_in <= 24'b100000101010000011010111;
#10000;
data_in <= 24'b011110011001100011001101;
#10000;
data_in <= 24'b011100001000111111000100;
#10000;
data_in <= 24'b011010001000011110111010;
#10000;
data_in <= 24'b011000101000000110110100;
#10000;
data_in <= 24'b010111010111110110101110;
#10000;
data_in <= 24'b010111000111101010101001;
#10000;
data_in <= 24'b100001101010010011011011;
#10000;
data_in <= 24'b100000001001111011010101;
#10000;
data_in <= 24'b011110001001011011001101;
#10000;
data_in <= 24'b011011111000111011000011;
#10000;
data_in <= 24'b011001111000100010111010;
#10000;
data_in <= 24'b011000011000001010110100;
#10000;
data_in <= 24'b010111010111111010101111;
#10000;
data_in <= 24'b010110110111110010101010;
#10000;
data_in <= 24'b100001001010001011011001;
#10000;
data_in <= 24'b011111111001110111010100;
#10000;
data_in <= 24'b011101111001010111001100;
#10000;
data_in <= 24'b011011111000111011000011;
#10000;
data_in <= 24'b011010001000100010111101;
#10000;
data_in <= 24'b011000111000010010110110;
#10000;
data_in <= 24'b010111111000000010110001;
#10000;
data_in <= 24'b010111100111111010101111;
#10000;
data_in <= 24'b100000111010000111011000;
#10000;
data_in <= 24'b011111101001101111010100;
#10000;
data_in <= 24'b011101101001010011001011;
#10000;
data_in <= 24'b011011111000111011000011;
#10000;
data_in <= 24'b011010011000100110111110;
#10000;
data_in <= 24'b011001001000010110110111;
#10000;
data_in <= 24'b010111111000001110110011;
#10000;
data_in <= 24'b010111111000000010110001;
#10000;
data_in <= 24'b100000101010000011010111;
#10000;
data_in <= 24'b011111011001101111010010;
#10000;
data_in <= 24'b011101101001010011001011;
#10000;
data_in <= 24'b011011101000111011000011;
#10000;
data_in <= 24'b011010011000101010111100;
#10000;
data_in <= 24'b011001001000011110111001;
#10000;
data_in <= 24'b011000011000010110110101;
#10000;
data_in <= 24'b011000011000001010110011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010111000111010110011111;
#10000;
data_in <= 24'b010110000111000010011010;
#10000;
data_in <= 24'b010011010110011010010000;
#10000;
data_in <= 24'b010011010110100010010100;
#10000;
data_in <= 24'b010110110111100010100100;
#10000;
data_in <= 24'b010111111000000110101100;
#10000;
data_in <= 24'b011000101000010010101111;
#10000;
data_in <= 24'b011010011000110010110111;
#10000;
data_in <= 24'b011000000111100110100101;
#10000;
data_in <= 24'b010110010111001010011110;
#10000;
data_in <= 24'b010010100110010110010001;
#10000;
data_in <= 24'b010010010110010010010000;
#10000;
data_in <= 24'b010101010111001010011110;
#10000;
data_in <= 24'b011000001000000010101011;
#10000;
data_in <= 24'b011010111000110110111000;
#10000;
data_in <= 24'b011110101001110111000101;
#10000;
data_in <= 24'b010111100111100010100110;
#10000;
data_in <= 24'b010110110111010010100000;
#10000;
data_in <= 24'b010011010110100010010100;
#10000;
data_in <= 24'b010010010110010010010000;
#10000;
data_in <= 24'b010100010110111010011010;
#10000;
data_in <= 24'b010111100111101110100111;
#10000;
data_in <= 24'b011011111000111110111000;
#10000;
data_in <= 24'b100001101010011111001110;
#10000;
data_in <= 24'b010111000111011010100100;
#10000;
data_in <= 24'b010111000111010010100010;
#10000;
data_in <= 24'b010100100110110110011001;
#10000;
data_in <= 24'b010011100110100110010101;
#10000;
data_in <= 24'b010100100110110110011001;
#10000;
data_in <= 24'b010110010111010110011110;
#10000;
data_in <= 24'b011011011000101010110001;
#10000;
data_in <= 24'b100010001010010111001010;
#10000;
data_in <= 24'b010110110111100010100101;
#10000;
data_in <= 24'b010111010111011110100101;
#10000;
data_in <= 24'b010101100111000110011101;
#10000;
data_in <= 24'b010100010110110010011000;
#10000;
data_in <= 24'b010100000110110010010101;
#10000;
data_in <= 24'b010101100111000010011000;
#10000;
data_in <= 24'b011011001000011110101100;
#10000;
data_in <= 24'b100011011010011111001011;
#10000;
data_in <= 24'b011000000111110010101011;
#10000;
data_in <= 24'b011000000111101010101000;
#10000;
data_in <= 24'b010110000111001110011111;
#10000;
data_in <= 24'b010100010110110110010110;
#10000;
data_in <= 24'b010100000110101010010010;
#10000;
data_in <= 24'b010101000110111010010011;
#10000;
data_in <= 24'b011011101000100010101100;
#10000;
data_in <= 24'b100101001010110111001111;
#10000;
data_in <= 24'b011000010111110110101100;
#10000;
data_in <= 24'b011000100111110010101010;
#10000;
data_in <= 24'b010111010111011010100010;
#10000;
data_in <= 24'b010101110111000010011010;
#10000;
data_in <= 24'b010100110110110010010100;
#10000;
data_in <= 24'b010100100110110010010001;
#10000;
data_in <= 24'b011010101000001110100101;
#10000;
data_in <= 24'b100011111010011011000110;
#10000;
data_in <= 24'b010111010111101110101010;
#10000;
data_in <= 24'b011000000111110010101011;
#10000;
data_in <= 24'b010111100111100010100110;
#10000;
data_in <= 24'b010110110111011010100010;
#10000;
data_in <= 24'b010101100111000010011000;
#10000;
data_in <= 24'b010011110110100110001110;
#10000;
data_in <= 24'b010111110111100010011010;
#10000;
data_in <= 24'b100000001001011110110111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011101111001100111000100;
#10000;
data_in <= 24'b100000001010001011001101;
#10000;
data_in <= 24'b011110011001100111000010;
#10000;
data_in <= 24'b011101111001011010111101;
#10000;
data_in <= 24'b100011011010101011001111;
#10000;
data_in <= 24'b011010011000010010101001;
#10000;
data_in <= 24'b000111010011010101011001;
#10000;
data_in <= 24'b000010010010000101000101;
#10000;
data_in <= 24'b100010111010101111010100;
#10000;
data_in <= 24'b100001111010011111010000;
#10000;
data_in <= 24'b100010011010100011001111;
#10000;
data_in <= 24'b100010011010011011001011;
#10000;
data_in <= 24'b100100011010110011010001;
#10000;
data_in <= 24'b011110011001001110110111;
#10000;
data_in <= 24'b001110110101001101110111;
#10000;
data_in <= 24'b000110010010111101010010;
#10000;
data_in <= 24'b100101001011001111011010;
#10000;
data_in <= 24'b100100011010111011010011;
#10000;
data_in <= 24'b100111111011101111011110;
#10000;
data_in <= 24'b100111101011100111011011;
#10000;
data_in <= 24'b100110001011000111010011;
#10000;
data_in <= 24'b100001101001110110111101;
#10000;
data_in <= 24'b010011000110000110000001;
#10000;
data_in <= 24'b000101110010110001001100;
#10000;
data_in <= 24'b100101111011001111010110;
#10000;
data_in <= 24'b101001011100000111100011;
#10000;
data_in <= 24'b101101111101000011110010;
#10000;
data_in <= 24'b101011011100010011100100;
#10000;
data_in <= 24'b101000011011011011010101;
#10000;
data_in <= 24'b100000111001011110110110;
#10000;
data_in <= 24'b001111000100111001101011;
#10000;
data_in <= 24'b000001100001100000110101;
#10000;
data_in <= 24'b101000001011100111011011;
#10000;
data_in <= 24'b110000001101101011111000;
#10000;
data_in <= 24'b110001001101100111111000;
#10000;
data_in <= 24'b101001011011101011010110;
#10000;
data_in <= 24'b100110011010110011000111;
#10000;
data_in <= 24'b011011111000000010011011;
#10000;
data_in <= 24'b001000000010111101001001;
#10000;
data_in <= 24'b000000000000110100100111;
#10000;
data_in <= 24'b101010001100000011011110;
#10000;
data_in <= 24'b110000011101011111110011;
#10000;
data_in <= 24'b101010011011111011011001;
#10000;
data_in <= 24'b011110001000110010100101;
#10000;
data_in <= 24'b011011100111110110010111;
#10000;
data_in <= 24'b010010010101011101101110;
#10000;
data_in <= 24'b000010000001010000101100;
#10000;
data_in <= 24'b000000000000100100011111;
#10000;
data_in <= 24'b101001001011101011010110;
#10000;
data_in <= 24'b100111001011000111001100;
#10000;
data_in <= 24'b011101111000100110100000;
#10000;
data_in <= 24'b001111110101000001100101;
#10000;
data_in <= 24'b001011010011101001010000;
#10000;
data_in <= 24'b000111100010100100111101;
#10000;
data_in <= 24'b000000000000100000011100;
#10000;
data_in <= 24'b000000000000010100011001;
#10000;
data_in <= 24'b100111011011001011001110;
#10000;
data_in <= 24'b011110001000110010100101;
#10000;
data_in <= 24'b010100000110000101110110;
#10000;
data_in <= 24'b000111000010101000111101;
#10000;
data_in <= 24'b000000100000111000100000;
#10000;
data_in <= 24'b000010000001000000100001;
#10000;
data_in <= 24'b000000010000100000011001;
#10000;
data_in <= 24'b000000000000001100010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000011010001110000101100;
#10000;
data_in <= 24'b000100110010001000110010;
#10000;
data_in <= 24'b001000100011001001000011;
#10000;
data_in <= 24'b001011010011110001001111;
#10000;
data_in <= 24'b000111110011000001000101;
#10000;
data_in <= 24'b000011100010000000110111;
#10000;
data_in <= 24'b000101100010101001000011;
#10000;
data_in <= 24'b001011000100000101011100;
#10000;
data_in <= 24'b000100100001111100101101;
#10000;
data_in <= 24'b000101000010000100101111;
#10000;
data_in <= 24'b000111100010110100111101;
#10000;
data_in <= 24'b001010100011100101001001;
#10000;
data_in <= 24'b001000100011000101000100;
#10000;
data_in <= 24'b000100110010001000110101;
#10000;
data_in <= 24'b000101000010010000111011;
#10000;
data_in <= 24'b001000100011001101001101;
#10000;
data_in <= 24'b000101010010001000110000;
#10000;
data_in <= 24'b000100100001111100101101;
#10000;
data_in <= 24'b000110100010011100110111;
#10000;
data_in <= 24'b001001100011010101000101;
#10000;
data_in <= 24'b001000110011001001000101;
#10000;
data_in <= 24'b000101000010001100110110;
#10000;
data_in <= 24'b000011010001110100110100;
#10000;
data_in <= 24'b000100010010001000111100;
#10000;
data_in <= 24'b000101000010000100101111;
#10000;
data_in <= 24'b000100000001110100101011;
#10000;
data_in <= 24'b000101110010010000110100;
#10000;
data_in <= 24'b001001010011001001000010;
#10000;
data_in <= 24'b001001000011001001000100;
#10000;
data_in <= 24'b000101010010010000110111;
#10000;
data_in <= 24'b000010110001100100101111;
#10000;
data_in <= 24'b000010100001101000110001;
#10000;
data_in <= 24'b000100010001111000101100;
#10000;
data_in <= 24'b000011110001110000101010;
#10000;
data_in <= 24'b000101100010001100110011;
#10000;
data_in <= 24'b001000110011000001000000;
#10000;
data_in <= 24'b001000100011000001000010;
#10000;
data_in <= 24'b000101010010010000110111;
#10000;
data_in <= 24'b000011010001110000101111;
#10000;
data_in <= 24'b000010110001110000110001;
#10000;
data_in <= 24'b000100010001111000101100;
#10000;
data_in <= 24'b000011100001101100101001;
#10000;
data_in <= 24'b000101000010000100110001;
#10000;
data_in <= 24'b000111100010101100111011;
#10000;
data_in <= 24'b001000010010110100111111;
#10000;
data_in <= 24'b000101110010010100110111;
#10000;
data_in <= 24'b000100010001111100110010;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b000101010010001000110010;
#10000;
data_in <= 24'b000011100001101100101011;
#10000;
data_in <= 24'b000100010001101100101100;
#10000;
data_in <= 24'b000110100010010000110101;
#10000;
data_in <= 24'b001000000010101000111011;
#10000;
data_in <= 24'b000110110010100000111000;
#10000;
data_in <= 24'b000101100010001000110100;
#10000;
data_in <= 24'b000100110010000100110100;
#10000;
data_in <= 24'b000110000010010100110101;
#10000;
data_in <= 24'b000011100001101100101011;
#10000;
data_in <= 24'b000011000001011000100111;
#10000;
data_in <= 24'b000101010001111100110000;
#10000;
data_in <= 24'b000111100010100000111001;
#10000;
data_in <= 24'b000111100010100000111001;
#10000;
data_in <= 24'b000110010010001100110100;
#10000;
data_in <= 24'b000101000010000000110010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010101000110100010000111;
#10000;
data_in <= 24'b010111000111000110010000;
#10000;
data_in <= 24'b010110010110111010001110;
#10000;
data_in <= 24'b010010010101111001111110;
#10000;
data_in <= 24'b001111110101010001110100;
#10000;
data_in <= 24'b010000010101011001110110;
#10000;
data_in <= 24'b010000000101010101110101;
#10000;
data_in <= 24'b001111000100111001101011;
#10000;
data_in <= 24'b010010000101101101110110;
#10000;
data_in <= 24'b010110010110101110001000;
#10000;
data_in <= 24'b010110100110111010001101;
#10000;
data_in <= 24'b010010010101110101111100;
#10000;
data_in <= 24'b001111110101010001110100;
#10000;
data_in <= 24'b010000110101100001111000;
#10000;
data_in <= 24'b010000010101010101111000;
#10000;
data_in <= 24'b001110000100101001101001;
#10000;
data_in <= 24'b001100010100010001011111;
#10000;
data_in <= 24'b010100000110001001111111;
#10000;
data_in <= 24'b010110110110111110001110;
#10000;
data_in <= 24'b010010110101111101111110;
#10000;
data_in <= 24'b001111100101001101110011;
#10000;
data_in <= 24'b010001000101100101111001;
#10000;
data_in <= 24'b010000010101011001110110;
#10000;
data_in <= 24'b001101000100011001100011;
#10000;
data_in <= 24'b000110110010110001000110;
#10000;
data_in <= 24'b010001000101011101110010;
#10000;
data_in <= 24'b010111110111000110001110;
#10000;
data_in <= 24'b010011110110001110000010;
#10000;
data_in <= 24'b010000000101010001110011;
#10000;
data_in <= 24'b010000010101011001110110;
#10000;
data_in <= 24'b001111100101001101110011;
#10000;
data_in <= 24'b001100100100011101100011;
#10000;
data_in <= 24'b000010110001101100110010;
#10000;
data_in <= 24'b001101110100100001100010;
#10000;
data_in <= 24'b010110010110110010000111;
#10000;
data_in <= 24'b010100110110100010000100;
#10000;
data_in <= 24'b010000100101011001110101;
#10000;
data_in <= 24'b001111010101000101110000;
#10000;
data_in <= 24'b001110100100111101101111;
#10000;
data_in <= 24'b001101100100101101100111;
#10000;
data_in <= 24'b000000100001000000100110;
#10000;
data_in <= 24'b001001000011010001001011;
#10000;
data_in <= 24'b010010100101101101110101;
#10000;
data_in <= 24'b010101010110100010000011;
#10000;
data_in <= 24'b010010000101110101111001;
#10000;
data_in <= 24'b001110110100111101101110;
#10000;
data_in <= 24'b001101110100110001101100;
#10000;
data_in <= 24'b001110110101000001101100;
#10000;
data_in <= 24'b000000000000110100100000;
#10000;
data_in <= 24'b000011100001111100110100;
#10000;
data_in <= 24'b001100010100001001011100;
#10000;
data_in <= 24'b010100000110001101111110;
#10000;
data_in <= 24'b010100000110010110000001;
#10000;
data_in <= 24'b001111000101000101101101;
#10000;
data_in <= 24'b001101000100100101101000;
#10000;
data_in <= 24'b001111100101001101101111;
#10000;
data_in <= 24'b000000000000110100011111;
#10000;
data_in <= 24'b000000010001000000100011;
#10000;
data_in <= 24'b001000000011000001000111;
#10000;
data_in <= 24'b010011010101111001111000;
#10000;
data_in <= 24'b010101110110101010000101;
#10000;
data_in <= 24'b001111100101001101101111;
#10000;
data_in <= 24'b001100110100100001100111;
#10000;
data_in <= 24'b010000000101010101110001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001110110100100101100000;
#10000;
data_in <= 24'b001011000011100001001010;
#10000;
data_in <= 24'b001000000010101000111011;
#10000;
data_in <= 24'b001001110011000000111110;
#10000;
data_in <= 24'b001101000011110101000111;
#10000;
data_in <= 24'b001101110100000101001000;
#10000;
data_in <= 24'b001100000011100000111111;
#10000;
data_in <= 24'b001001100010111000110101;
#10000;
data_in <= 24'b001100010011111101010101;
#10000;
data_in <= 24'b001010110011011101001001;
#10000;
data_in <= 24'b001010000011001001000011;
#10000;
data_in <= 24'b001011010011011001000011;
#10000;
data_in <= 24'b001011110011100001000001;
#10000;
data_in <= 24'b001001110010111100110110;
#10000;
data_in <= 24'b000101110001110100100010;
#10000;
data_in <= 24'b000010000001000100010101;
#10000;
data_in <= 24'b001011110011110101010100;
#10000;
data_in <= 24'b001011000011100001001010;
#10000;
data_in <= 24'b001010010011001101000100;
#10000;
data_in <= 24'b001001100010111100111100;
#10000;
data_in <= 24'b000111100010011100110001;
#10000;
data_in <= 24'b000100100001110000100011;
#10000;
data_in <= 24'b000010110001001100011010;
#10000;
data_in <= 24'b000010000001000000010111;
#10000;
data_in <= 24'b001100000100000001010111;
#10000;
data_in <= 24'b001011110011110101010000;
#10000;
data_in <= 24'b001010010011011001000110;
#10000;
data_in <= 24'b000111100010100100110111;
#10000;
data_in <= 24'b000100000001101000100100;
#10000;
data_in <= 24'b000001110001000000011001;
#10000;
data_in <= 24'b000010010001001000011011;
#10000;
data_in <= 24'b000100100001101100100100;
#10000;
data_in <= 24'b001100110100001101011010;
#10000;
data_in <= 24'b001101000100001001010101;
#10000;
data_in <= 24'b001011010011101101001101;
#10000;
data_in <= 24'b000111110010110000111100;
#10000;
data_in <= 24'b000011000001011100100101;
#10000;
data_in <= 24'b000000000000100100010110;
#10000;
data_in <= 24'b000000100000101100011000;
#10000;
data_in <= 24'b000010010001010100100001;
#10000;
data_in <= 24'b001110010100100001100010;
#10000;
data_in <= 24'b001100110100000101010111;
#10000;
data_in <= 24'b001010000011011001001001;
#10000;
data_in <= 24'b000101110010010100110111;
#10000;
data_in <= 24'b000001110001010000100100;
#10000;
data_in <= 24'b000000000000110100011101;
#10000;
data_in <= 24'b000001110001010000100010;
#10000;
data_in <= 24'b000100110010000000101110;
#10000;
data_in <= 24'b001111100100111101101001;
#10000;
data_in <= 24'b001101000100010101011010;
#10000;
data_in <= 24'b001001110011010101001011;
#10000;
data_in <= 24'b000110100010100100111100;
#10000;
data_in <= 24'b000100110010000100110100;
#10000;
data_in <= 24'b000101000010001000110100;
#10000;
data_in <= 24'b000111100010110000111110;
#10000;
data_in <= 24'b001010010011100101001010;
#10000;
data_in <= 24'b010000000101000101101011;
#10000;
data_in <= 24'b001110110100101101100010;
#10000;
data_in <= 24'b001101000100010001011011;
#10000;
data_in <= 24'b001100000100000001010111;
#10000;
data_in <= 24'b001011010011111001010011;
#10000;
data_in <= 24'b001010100011101101010000;
#10000;
data_in <= 24'b001010010011101001001111;
#10000;
data_in <= 24'b001010110011101101010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000011010001011000011111;
#10000;
data_in <= 24'b000001000000111000011000;
#10000;
data_in <= 24'b000000000000001000010011;
#10000;
data_in <= 24'b000000000000011100011010;
#10000;
data_in <= 24'b000101110010011001000000;
#10000;
data_in <= 24'b010010000101011101110111;
#10000;
data_in <= 24'b011011010111110110100001;
#10000;
data_in <= 24'b011110101000111110101111;
#10000;
data_in <= 24'b000001010000111000010111;
#10000;
data_in <= 24'b000000000000011000010000;
#10000;
data_in <= 24'b000000000000101000011011;
#10000;
data_in <= 24'b000111000010100100111111;
#10000;
data_in <= 24'b010000010101001001101101;
#10000;
data_in <= 24'b010111110111001010010011;
#10000;
data_in <= 24'b011101011000100010101101;
#10000;
data_in <= 24'b100000001001011010111001;
#10000;
data_in <= 24'b000001110001000000011001;
#10000;
data_in <= 24'b000000010000110100011001;
#10000;
data_in <= 24'b000101010010000100110011;
#10000;
data_in <= 24'b001111110100110101100011;
#10000;
data_in <= 24'b010111000110110110001000;
#10000;
data_in <= 24'b011001100111100110011010;
#10000;
data_in <= 24'b011101001000011110101100;
#10000;
data_in <= 24'b100001001001110110111111;
#10000;
data_in <= 24'b000100100001110000100110;
#10000;
data_in <= 24'b000101110010001000110000;
#10000;
data_in <= 24'b001011010011101101001101;
#10000;
data_in <= 24'b010010110101101101110010;
#10000;
data_in <= 24'b010110100110101010000111;
#10000;
data_in <= 24'b011000000111001110010100;
#10000;
data_in <= 24'b011110101001000010110100;
#10000;
data_in <= 24'b100110011011000111010101;
#10000;
data_in <= 24'b000110000010001100110001;
#10000;
data_in <= 24'b001001000011000101000001;
#10000;
data_in <= 24'b001101110100011001011001;
#10000;
data_in <= 24'b010010010101101001110100;
#10000;
data_in <= 24'b010110110110110110001010;
#10000;
data_in <= 24'b011100111000011110101010;
#10000;
data_in <= 24'b100110001010111011010010;
#10000;
data_in <= 24'b101100111100110111110001;
#10000;
data_in <= 24'b001000010010110100111111;
#10000;
data_in <= 24'b001010110011101001001101;
#10000;
data_in <= 24'b001111000100110001100011;
#10000;
data_in <= 24'b010100000110001101111110;
#10000;
data_in <= 24'b011011111000010010100011;
#10000;
data_in <= 24'b100101001010101011001101;
#10000;
data_in <= 24'b101011011100010111101001;
#10000;
data_in <= 24'b101101011101000111110100;
#10000;
data_in <= 24'b001011010011101101010001;
#10000;
data_in <= 24'b001110010100100101100000;
#10000;
data_in <= 24'b010100000110000101111011;
#10000;
data_in <= 24'b011011001000000110011101;
#10000;
data_in <= 24'b100011111010011011000110;
#10000;
data_in <= 24'b101011001100010111100111;
#10000;
data_in <= 24'b101101111100111111110011;
#10000;
data_in <= 24'b101100011100110111110000;
#10000;
data_in <= 24'b001100100100001101011101;
#10000;
data_in <= 24'b010001010101100001110011;
#10000;
data_in <= 24'b011001100111101110010111;
#10000;
data_in <= 24'b100011001010000111000000;
#10000;
data_in <= 24'b101010001100000111100011;
#10000;
data_in <= 24'b101110011101001111110111;
#10000;
data_in <= 24'b101111101101100011111101;
#10000;
data_in <= 24'b101110011101011111111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100010011010000110111101;
#10000;
data_in <= 24'b100110111011100011010011;
#10000;
data_in <= 24'b101011001100101011100111;
#10000;
data_in <= 24'b101001101100011111101000;
#10000;
data_in <= 24'b100111001011111111100001;
#10000;
data_in <= 24'b100101001011100111011111;
#10000;
data_in <= 24'b100011101011010111011100;
#10000;
data_in <= 24'b100001111010111111011001;
#10000;
data_in <= 24'b100101101011000111001100;
#10000;
data_in <= 24'b101001001100001111011100;
#10000;
data_in <= 24'b101011101100111111101001;
#10000;
data_in <= 24'b101010001100101011101000;
#10000;
data_in <= 24'b100111001100000111100011;
#10000;
data_in <= 24'b100101001011101111100001;
#10000;
data_in <= 24'b100011111011011011011101;
#10000;
data_in <= 24'b100001111010111111011001;
#10000;
data_in <= 24'b101001111100010011011111;
#10000;
data_in <= 24'b101011111100111011100111;
#10000;
data_in <= 24'b101100011101001011101100;
#10000;
data_in <= 24'b101001111100101111101001;
#10000;
data_in <= 24'b100111101100001111100101;
#10000;
data_in <= 24'b100101101011110111100011;
#10000;
data_in <= 24'b100100001011011111011110;
#10000;
data_in <= 24'b100001101010111011011000;
#10000;
data_in <= 24'b101100111101000111101110;
#10000;
data_in <= 24'b101100111101010011101110;
#10000;
data_in <= 24'b101011101101000011101101;
#10000;
data_in <= 24'b101001101100101011101000;
#10000;
data_in <= 24'b100111101100010011100110;
#10000;
data_in <= 24'b100110001011111111100101;
#10000;
data_in <= 24'b100011101011011111011110;
#10000;
data_in <= 24'b100001101010111011011000;
#10000;
data_in <= 24'b101101011101010111110010;
#10000;
data_in <= 24'b101011111101010011101110;
#10000;
data_in <= 24'b101010011100111011101010;
#10000;
data_in <= 24'b101000101100100011101000;
#10000;
data_in <= 24'b100111111100010111100111;
#10000;
data_in <= 24'b100110011100000011100110;
#10000;
data_in <= 24'b100011101011011111011110;
#10000;
data_in <= 24'b100001011010110111010111;
#10000;
data_in <= 24'b101100101101010011110001;
#10000;
data_in <= 24'b101010101101000111101101;
#10000;
data_in <= 24'b101001101100110011101010;
#10000;
data_in <= 24'b101000111100101011101010;
#10000;
data_in <= 24'b100111111100100011101001;
#10000;
data_in <= 24'b100110101100000111100111;
#10000;
data_in <= 24'b100011101011011111011110;
#10000;
data_in <= 24'b100001011010110111010111;
#10000;
data_in <= 24'b101011111101001111110001;
#10000;
data_in <= 24'b101010011101000111101101;
#10000;
data_in <= 24'b101001111100111111101100;
#10000;
data_in <= 24'b101001011100111011101110;
#10000;
data_in <= 24'b101001001100110111101110;
#10000;
data_in <= 24'b100111011100010011101010;
#10000;
data_in <= 24'b100100011011100011011111;
#10000;
data_in <= 24'b100010001010111111010110;
#10000;
data_in <= 24'b101011011101001111110001;
#10000;
data_in <= 24'b101010101101001011101111;
#10000;
data_in <= 24'b101010001101000111110001;
#10000;
data_in <= 24'b101010101101001111110100;
#10000;
data_in <= 24'b101010001101000011110011;
#10000;
data_in <= 24'b100111111100011111101010;
#10000;
data_in <= 24'b100100101011100111100000;
#10000;
data_in <= 24'b100010001010111111010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100001111010111011011010;
#10000;
data_in <= 24'b100011111011011011100010;
#10000;
data_in <= 24'b100101101011110011100110;
#10000;
data_in <= 24'b100111001100000011101000;
#10000;
data_in <= 24'b101010101100111011110100;
#10000;
data_in <= 24'b101110101101110011111111;
#10000;
data_in <= 24'b101110111101100111111100;
#10000;
data_in <= 24'b101011101100101111110000;
#10000;
data_in <= 24'b100000011010101111010110;
#10000;
data_in <= 24'b100010001010111111011011;
#10000;
data_in <= 24'b100100001011011011100000;
#10000;
data_in <= 24'b100110001011110011100100;
#10000;
data_in <= 24'b101001001100010111101100;
#10000;
data_in <= 24'b101011101100111011110010;
#10000;
data_in <= 24'b101100111101000111110100;
#10000;
data_in <= 24'b101100011100111011110011;
#10000;
data_in <= 24'b100001011010110011011000;
#10000;
data_in <= 24'b100010011011000011011100;
#10000;
data_in <= 24'b100100101011100011100010;
#10000;
data_in <= 24'b100111001100000011101000;
#10000;
data_in <= 24'b101000101100001111101010;
#10000;
data_in <= 24'b101001001100010011101000;
#10000;
data_in <= 24'b101001101100010011100111;
#10000;
data_in <= 24'b101001101100001111101000;
#10000;
data_in <= 24'b100010001010111111011011;
#10000;
data_in <= 24'b100011111011010011100000;
#10000;
data_in <= 24'b100101101011100111100100;
#10000;
data_in <= 24'b100110101011110111100101;
#10000;
data_in <= 24'b101000001011111111100110;
#10000;
data_in <= 24'b100111101011101111100000;
#10000;
data_in <= 24'b100100111010111011010011;
#10000;
data_in <= 24'b100001001010000111000110;
#10000;
data_in <= 24'b100010011010111011011010;
#10000;
data_in <= 24'b100010111011000011011100;
#10000;
data_in <= 24'b100010001010101111010110;
#10000;
data_in <= 24'b100001001010011111001111;
#10000;
data_in <= 24'b100010101010100111010000;
#10000;
data_in <= 24'b100011001010100111001110;
#10000;
data_in <= 24'b011111001001011110111100;
#10000;
data_in <= 24'b011001011000000010100101;
#10000;
data_in <= 24'b100010011010111011011010;
#10000;
data_in <= 24'b100001001010011111010011;
#10000;
data_in <= 24'b011101111001100111000100;
#10000;
data_in <= 24'b011010111000101110110110;
#10000;
data_in <= 24'b011011001000100010110001;
#10000;
data_in <= 24'b011011001000011010101110;
#10000;
data_in <= 24'b011000100111101110100011;
#10000;
data_in <= 24'b010100010110101110010011;
#10000;
data_in <= 24'b100010111010111011011001;
#10000;
data_in <= 24'b011111001001111111001010;
#10000;
data_in <= 24'b011011001000111010111001;
#10000;
data_in <= 24'b010111100111111010101001;
#10000;
data_in <= 24'b010011000110100010010001;
#10000;
data_in <= 24'b001110010101001101111011;
#10000;
data_in <= 24'b001101010100111001110110;
#10000;
data_in <= 24'b001111000101010101111101;
#10000;
data_in <= 24'b100010001010101111010110;
#10000;
data_in <= 24'b011101101001100011000011;
#10000;
data_in <= 24'b011010101000101010110101;
#10000;
data_in <= 24'b010111000111100110100101;
#10000;
data_in <= 24'b001101100101001001111011;
#10000;
data_in <= 24'b000010110010010001001110;
#10000;
data_in <= 24'b000010000010000001001010;
#10000;
data_in <= 24'b001000010011101001100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101010011100011011110010;
#10000;
data_in <= 24'b100101001011001111100000;
#10000;
data_in <= 24'b011110101001100111000110;
#10000;
data_in <= 24'b011010011000100010110101;
#10000;
data_in <= 24'b011011011000101110111010;
#10000;
data_in <= 24'b011110001001011011000101;
#10000;
data_in <= 24'b011111001001101011001001;
#10000;
data_in <= 24'b011110001001011111000100;
#10000;
data_in <= 24'b100111101011110011100101;
#10000;
data_in <= 24'b011101101001010111000010;
#10000;
data_in <= 24'b010101110111011010100011;
#10000;
data_in <= 24'b010101110111011010100011;
#10000;
data_in <= 24'b011000101000000010101111;
#10000;
data_in <= 24'b011010011000011110110110;
#10000;
data_in <= 24'b011100111000111110111110;
#10000;
data_in <= 24'b011111001001100011000111;
#10000;
data_in <= 24'b100011001010101011010011;
#10000;
data_in <= 24'b011010101000101010110101;
#10000;
data_in <= 24'b010010100110100110010110;
#10000;
data_in <= 24'b001111110101111010001011;
#10000;
data_in <= 24'b001111000101101010001001;
#10000;
data_in <= 24'b001111010101101110001010;
#10000;
data_in <= 24'b010010000110011010010101;
#10000;
data_in <= 24'b010101110111010110100100;
#10000;
data_in <= 24'b011010001000011010101111;
#10000;
data_in <= 24'b010111100111111010101001;
#10000;
data_in <= 24'b001111110101111010001011;
#10000;
data_in <= 24'b000100010011000001011101;
#10000;
data_in <= 24'b000000000001001101000010;
#10000;
data_in <= 24'b000000000001101001001001;
#10000;
data_in <= 24'b000110000011011001100101;
#10000;
data_in <= 24'b001011100100110001111011;
#10000;
data_in <= 24'b010101000111000010011001;
#10000;
data_in <= 24'b010100000110111010010111;
#10000;
data_in <= 24'b001100110101000001111100;
#10000;
data_in <= 24'b000000000001110101001001;
#10000;
data_in <= 24'b000000000000000000101000;
#10000;
data_in <= 24'b000000000000011100110100;
#10000;
data_in <= 24'b000011000010110101011011;
#10000;
data_in <= 24'b001010100100101101111001;
#10000;
data_in <= 24'b010010000110010110001100;
#10000;
data_in <= 24'b001110110101100110000010;
#10000;
data_in <= 24'b001010110100100001110100;
#10000;
data_in <= 24'b000101110011010001100000;
#10000;
data_in <= 24'b000000010010000001001101;
#10000;
data_in <= 24'b000000000001101101001000;
#10000;
data_in <= 24'b000010110010110001011010;
#10000;
data_in <= 24'b001000010100001101110001;
#10000;
data_in <= 24'b001101000101000101111000;
#10000;
data_in <= 24'b001010110100101001110001;
#10000;
data_in <= 24'b001001010100001101101100;
#10000;
data_in <= 24'b001000110100000001101100;
#10000;
data_in <= 24'b000111110011111001101011;
#10000;
data_in <= 24'b000111110011111001101011;
#10000;
data_in <= 24'b001001000100010101110011;
#10000;
data_in <= 24'b001011010100111101111101;
#10000;
data_in <= 24'b001100110101000001110111;
#10000;
data_in <= 24'b001101100101010101111100;
#10000;
data_in <= 24'b001011110100110101110110;
#10000;
data_in <= 24'b001001000100000101101101;
#10000;
data_in <= 24'b001011100100110101111010;
#10000;
data_in <= 24'b010011110111000010011110;
#10000;
data_in <= 24'b011011001000110110111011;
#10000;
data_in <= 24'b011101101001100011000110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011101111001011011000011;
#10000;
data_in <= 24'b100101011011001011011110;
#10000;
data_in <= 24'b101001011100001111101100;
#10000;
data_in <= 24'b101010001100010111101010;
#10000;
data_in <= 24'b101011011100101111101110;
#10000;
data_in <= 24'b101100111101001011110011;
#10000;
data_in <= 24'b101101001101001111110100;
#10000;
data_in <= 24'b101101001101001111110100;
#10000;
data_in <= 24'b011011011000101010110111;
#10000;
data_in <= 24'b100000001001110111001001;
#10000;
data_in <= 24'b100110011011011011100010;
#10000;
data_in <= 24'b101010001100011111101110;
#10000;
data_in <= 24'b101011011100101011110001;
#10000;
data_in <= 24'b101011001100110011110000;
#10000;
data_in <= 24'b101011101100110011101111;
#10000;
data_in <= 24'b101010101100101011101101;
#10000;
data_in <= 24'b010101010111010010100001;
#10000;
data_in <= 24'b010111000111110010100111;
#10000;
data_in <= 24'b100000001010000011001011;
#10000;
data_in <= 24'b101000111100010011101011;
#10000;
data_in <= 24'b101010111100101011110001;
#10000;
data_in <= 24'b101010001100101011101110;
#10000;
data_in <= 24'b101011111100111111110010;
#10000;
data_in <= 24'b101010111100111011110000;
#10000;
data_in <= 24'b010000010110000010001101;
#10000;
data_in <= 24'b001111010101111010001011;
#10000;
data_in <= 24'b011010101000110010110111;
#10000;
data_in <= 24'b100111011100000011101000;
#10000;
data_in <= 24'b101001011100100111101111;
#10000;
data_in <= 24'b101001101100101011101110;
#10000;
data_in <= 24'b101011111101001111110111;
#10000;
data_in <= 24'b101011101101001011110110;
#10000;
data_in <= 24'b001010110100110001111001;
#10000;
data_in <= 24'b001011010101000001111100;
#10000;
data_in <= 24'b011000011000010010101111;
#10000;
data_in <= 24'b100110101011111011100110;
#10000;
data_in <= 24'b101001001100100111101111;
#10000;
data_in <= 24'b101001001100101011101101;
#10000;
data_in <= 24'b101010111101000111110100;
#10000;
data_in <= 24'b101010001100111011110001;
#10000;
data_in <= 24'b001000100100010101110001;
#10000;
data_in <= 24'b001100000101010110000001;
#10000;
data_in <= 24'b011001001000100110110101;
#10000;
data_in <= 24'b100101111011110111100111;
#10000;
data_in <= 24'b101001011100110011110011;
#10000;
data_in <= 24'b101001011100111111110100;
#10000;
data_in <= 24'b101001111101000111110110;
#10000;
data_in <= 24'b101001001100101111110001;
#10000;
data_in <= 24'b010001100110100010010110;
#10000;
data_in <= 24'b010111011000001010101110;
#10000;
data_in <= 24'b100000001010010111010001;
#10000;
data_in <= 24'b100101111011111111101001;
#10000;
data_in <= 24'b101000011100100111110011;
#10000;
data_in <= 24'b101000111100111011110101;
#10000;
data_in <= 24'b101000101100110111110100;
#10000;
data_in <= 24'b100111111100101011110001;
#10000;
data_in <= 24'b011111101010001011010010;
#10000;
data_in <= 24'b100101101011101011101000;
#10000;
data_in <= 24'b101000001100011111110100;
#10000;
data_in <= 24'b100110111100001011101110;
#10000;
data_in <= 24'b100110011100001111101110;
#10000;
data_in <= 24'b100110111100010111110000;
#10000;
data_in <= 24'b100101111100001111101100;
#10000;
data_in <= 24'b100101101100001011101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101001111100011111101011;
#10000;
data_in <= 24'b101001101100010111101100;
#10000;
data_in <= 24'b101000101100001111101010;
#10000;
data_in <= 24'b100111111011111111101010;
#10000;
data_in <= 24'b100110111011101011100111;
#10000;
data_in <= 24'b100101101011010011100101;
#10000;
data_in <= 24'b100011011010110011011111;
#10000;
data_in <= 24'b100010011010100011011101;
#10000;
data_in <= 24'b101010101100100111110000;
#10000;
data_in <= 24'b101001101100011111101110;
#10000;
data_in <= 24'b101000111100001111101100;
#10000;
data_in <= 24'b100111111011111111101010;
#10000;
data_in <= 24'b100110111011101011100111;
#10000;
data_in <= 24'b100101011011001111100010;
#10000;
data_in <= 24'b100011011010110111011110;
#10000;
data_in <= 24'b100010011010100011011011;
#10000;
data_in <= 24'b101010101100101111110010;
#10000;
data_in <= 24'b101001011100100111101111;
#10000;
data_in <= 24'b101000001100001111101011;
#10000;
data_in <= 24'b100110111011110111101000;
#10000;
data_in <= 24'b100101101011011111100100;
#10000;
data_in <= 24'b100100001011000111011111;
#10000;
data_in <= 24'b100010111010101111011100;
#10000;
data_in <= 24'b100001111010011111011000;
#10000;
data_in <= 24'b101010011100110111110011;
#10000;
data_in <= 24'b101001011100100111101111;
#10000;
data_in <= 24'b100111111100001011101010;
#10000;
data_in <= 24'b100110001011101011100101;
#10000;
data_in <= 24'b100100111011010011100001;
#10000;
data_in <= 24'b100011101010111111011101;
#10000;
data_in <= 24'b100010011010100111011010;
#10000;
data_in <= 24'b100001101010011011010111;
#10000;
data_in <= 24'b101010101100111111110101;
#10000;
data_in <= 24'b101001011100100111110001;
#10000;
data_in <= 24'b100111101100000111101100;
#10000;
data_in <= 24'b100101111011101011100101;
#10000;
data_in <= 24'b100100101011010111100001;
#10000;
data_in <= 24'b100011011011000011011100;
#10000;
data_in <= 24'b100010011010101111011001;
#10000;
data_in <= 24'b100001101010100011010110;
#10000;
data_in <= 24'b101010001100111111110110;
#10000;
data_in <= 24'b101001101100101011110010;
#10000;
data_in <= 24'b100111111100001011101101;
#10000;
data_in <= 24'b100110011011110011100111;
#10000;
data_in <= 24'b100101001011011111100011;
#10000;
data_in <= 24'b100100001011001111011111;
#10000;
data_in <= 24'b100011001010111011011100;
#10000;
data_in <= 24'b100010011010101111011001;
#10000;
data_in <= 24'b101000101100101111110010;
#10000;
data_in <= 24'b101000011100011111110001;
#10000;
data_in <= 24'b100111001100000111101101;
#10000;
data_in <= 24'b100101111011110011101000;
#10000;
data_in <= 24'b100100101011011111100011;
#10000;
data_in <= 24'b100011101011001111011111;
#10000;
data_in <= 24'b100011001010111111011011;
#10000;
data_in <= 24'b100010011010110011011000;
#10000;
data_in <= 24'b100111011100010011110000;
#10000;
data_in <= 24'b100110101100000111101101;
#10000;
data_in <= 24'b100110001011110111101001;
#10000;
data_in <= 24'b100101001011100111100101;
#10000;
data_in <= 24'b100100001011010111100001;
#10000;
data_in <= 24'b100011001011000111011101;
#10000;
data_in <= 24'b100010101010110111011001;
#10000;
data_in <= 24'b100001111010101011010110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100000001001111111010100;
#10000;
data_in <= 24'b011110111001101111010000;
#10000;
data_in <= 24'b011101011001010111001010;
#10000;
data_in <= 24'b011011011000111111000100;
#10000;
data_in <= 24'b011010001000101110111101;
#10000;
data_in <= 24'b011001001000011110111001;
#10000;
data_in <= 24'b011000001000010010110100;
#10000;
data_in <= 24'b010111101000001010110010;
#10000;
data_in <= 24'b100000001010000011010101;
#10000;
data_in <= 24'b011111001001110011010001;
#10000;
data_in <= 24'b011100111001010111001010;
#10000;
data_in <= 24'b011011011001000011000010;
#10000;
data_in <= 24'b011010001000101110111101;
#10000;
data_in <= 24'b011001001000100010111000;
#10000;
data_in <= 24'b011000011000010110110101;
#10000;
data_in <= 24'b010111111000001110110011;
#10000;
data_in <= 24'b100000011010001011010100;
#10000;
data_in <= 24'b011111001001110111001111;
#10000;
data_in <= 24'b011101001001010111000111;
#10000;
data_in <= 24'b011011101000111111000001;
#10000;
data_in <= 24'b011010011000101010111100;
#10000;
data_in <= 24'b011001101000011110111000;
#10000;
data_in <= 24'b011001001000010110110110;
#10000;
data_in <= 24'b011000101000010010110010;
#10000;
data_in <= 24'b100000101010001111010100;
#10000;
data_in <= 24'b011111001001110111001110;
#10000;
data_in <= 24'b011101001001010111000111;
#10000;
data_in <= 24'b011011011000111010111111;
#10000;
data_in <= 24'b011010011000101010111011;
#10000;
data_in <= 24'b011001101000100010110110;
#10000;
data_in <= 24'b011001011000011110110101;
#10000;
data_in <= 24'b011001001000011010110100;
#10000;
data_in <= 24'b100000111010010011010010;
#10000;
data_in <= 24'b011111011001111011001100;
#10000;
data_in <= 24'b011101011001010111000110;
#10000;
data_in <= 24'b011011101000111110111101;
#10000;
data_in <= 24'b011010101000101110111001;
#10000;
data_in <= 24'b011010001000100110110110;
#10000;
data_in <= 24'b011001101000011110110100;
#10000;
data_in <= 24'b011001011000011110110101;
#10000;
data_in <= 24'b100000101010001111010001;
#10000;
data_in <= 24'b011111011001111011001100;
#10000;
data_in <= 24'b011101101001011111000101;
#10000;
data_in <= 24'b011011111001000010111101;
#10000;
data_in <= 24'b011010111000110010111001;
#10000;
data_in <= 24'b011010011000101010110111;
#10000;
data_in <= 24'b011001111000100010110101;
#10000;
data_in <= 24'b011001101000011110110100;
#10000;
data_in <= 24'b100000011010001011001111;
#10000;
data_in <= 24'b011111001001110111001010;
#10000;
data_in <= 24'b011110001001011111000100;
#10000;
data_in <= 24'b011100111001001110111110;
#10000;
data_in <= 24'b011011111000111110111010;
#10000;
data_in <= 24'b011011001000110010110111;
#10000;
data_in <= 24'b011010011000100110110100;
#10000;
data_in <= 24'b011001111000011010110011;
#10000;
data_in <= 24'b100000001010000111001110;
#10000;
data_in <= 24'b011111001001110111001010;
#10000;
data_in <= 24'b011110001001100011000011;
#10000;
data_in <= 24'b011100111001001110111110;
#10000;
data_in <= 24'b011100001001000010111011;
#10000;
data_in <= 24'b011011001000110010110111;
#10000;
data_in <= 24'b011010111000100110110010;
#10000;
data_in <= 24'b011001111000011110110010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010110100111110010101010;
#10000;
data_in <= 24'b010111000111110110101011;
#10000;
data_in <= 24'b011000011000000010101101;
#10000;
data_in <= 24'b010111110111111110101010;
#10000;
data_in <= 24'b010110000111011010011111;
#10000;
data_in <= 24'b010100100110111110010110;
#10000;
data_in <= 24'b010110000111001010010110;
#10000;
data_in <= 24'b011001000111101010011101;
#10000;
data_in <= 24'b011000001000001010110000;
#10000;
data_in <= 24'b010111010111111110101101;
#10000;
data_in <= 24'b010111000111110110101011;
#10000;
data_in <= 24'b010110110111110010101001;
#10000;
data_in <= 24'b010110100111011110100011;
#10000;
data_in <= 24'b010100110111000010010111;
#10000;
data_in <= 24'b010100100110110110010010;
#10000;
data_in <= 24'b010101110111000010010010;
#10000;
data_in <= 24'b011000111000010010110101;
#10000;
data_in <= 24'b010111010111111110101101;
#10000;
data_in <= 24'b010110010111101010101000;
#10000;
data_in <= 24'b010110010111101010100111;
#10000;
data_in <= 24'b010111000111100110100101;
#10000;
data_in <= 24'b010110000111010010011101;
#10000;
data_in <= 24'b010100010110110010010001;
#10000;
data_in <= 24'b010011110110100010001010;
#10000;
data_in <= 24'b010111111000000010110001;
#10000;
data_in <= 24'b010110100111101110101100;
#10000;
data_in <= 24'b010110000111100010101001;
#10000;
data_in <= 24'b010110100111101110101001;
#10000;
data_in <= 24'b010111010111110010101001;
#10000;
data_in <= 24'b010111010111100110100010;
#10000;
data_in <= 24'b010101100111000110010110;
#10000;
data_in <= 24'b010100010110101010001100;
#10000;
data_in <= 24'b010111000111110110101110;
#10000;
data_in <= 24'b010110100111111010101110;
#10000;
data_in <= 24'b010111000111110110101110;
#10000;
data_in <= 24'b010111010111111010101100;
#10000;
data_in <= 24'b010111110111111010101011;
#10000;
data_in <= 24'b010111010111101110100100;
#10000;
data_in <= 24'b010110100111010110011010;
#10000;
data_in <= 24'b010101110111000010010010;
#10000;
data_in <= 24'b010111111000000010110001;
#10000;
data_in <= 24'b011000001000001110110101;
#10000;
data_in <= 24'b011000101000001110110101;
#10000;
data_in <= 24'b010111111000000110101111;
#10000;
data_in <= 24'b010111100111110110101010;
#10000;
data_in <= 24'b010111010111101110100100;
#10000;
data_in <= 24'b010110110111011010011011;
#10000;
data_in <= 24'b010110000111000110010001;
#10000;
data_in <= 24'b011000111000010010110101;
#10000;
data_in <= 24'b011000101000010110110111;
#10000;
data_in <= 24'b011000111000010010110110;
#10000;
data_in <= 24'b010111111000000010110001;
#10000;
data_in <= 24'b010111110111110110101100;
#10000;
data_in <= 24'b010111100111101110100111;
#10000;
data_in <= 24'b010110110111011010011011;
#10000;
data_in <= 24'b010101110111000010010000;
#10000;
data_in <= 24'b011000111000010010110110;
#10000;
data_in <= 24'b011000011000001110111000;
#10000;
data_in <= 24'b011000001000000110110011;
#10000;
data_in <= 24'b010111000111110110101110;
#10000;
data_in <= 24'b010111010111111010101100;
#10000;
data_in <= 24'b011000010111111110101000;
#10000;
data_in <= 24'b010111010111100010011101;
#10000;
data_in <= 24'b010101110111000010010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011011111000001110100010;
#10000;
data_in <= 24'b010111110111000010001010;
#10000;
data_in <= 24'b010001000101001001101000;
#10000;
data_in <= 24'b000110010010010100110111;
#10000;
data_in <= 24'b000000000000000000001111;
#10000;
data_in <= 24'b000000000000010100010010;
#10000;
data_in <= 24'b000010100000111100011000;
#10000;
data_in <= 24'b000000000000000000001001;
#10000;
data_in <= 24'b001111110101001101110010;
#10000;
data_in <= 24'b001001110011100001010010;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
data_in <= 24'b000010110001010100100110;
#10000;
data_in <= 24'b000000000000010000010001;
#10000;
data_in <= 24'b000000000000010100001110;
#10000;
data_in <= 24'b000010100000110000010100;
#10000;
data_in <= 24'b000001100000100100001110;
#10000;
data_in <= 24'b001101000100100101100101;
#10000;
data_in <= 24'b000010110001110000110110;
#10000;
data_in <= 24'b000000000000011100011010;
#10000;
data_in <= 24'b000000100000110000011101;
#10000;
data_in <= 24'b000001000000101000010101;
#10000;
data_in <= 24'b000000000000010000001011;
#10000;
data_in <= 24'b000000110000011000001011;
#10000;
data_in <= 24'b000010100000110100010001;
#10000;
data_in <= 24'b010011100110001101111111;
#10000;
data_in <= 24'b000110110010110101000100;
#10000;
data_in <= 24'b000000000000011100011010;
#10000;
data_in <= 24'b000000000000101000011000;
#10000;
data_in <= 24'b000001110000110100011000;
#10000;
data_in <= 24'b000000010000010000001100;
#10000;
data_in <= 24'b000000010000010000001000;
#10000;
data_in <= 24'b000010110000111100010000;
#10000;
data_in <= 24'b010110000110110110001001;
#10000;
data_in <= 24'b001010110011110101010100;
#10000;
data_in <= 24'b000000010000111100100001;
#10000;
data_in <= 24'b000000000000011100010011;
#10000;
data_in <= 24'b000001100000110100010110;
#10000;
data_in <= 24'b000001110000101100010000;
#10000;
data_in <= 24'b000001010000100100001010;
#10000;
data_in <= 24'b000011000000111000001110;
#10000;
data_in <= 24'b010100110110100010000100;
#10000;
data_in <= 24'b001101100100100101011110;
#10000;
data_in <= 24'b000011100001110100101101;
#10000;
data_in <= 24'b000000000000100000010010;
#10000;
data_in <= 24'b000001110000111100010110;
#10000;
data_in <= 24'b000011000001000100010100;
#10000;
data_in <= 24'b000010000000101000001010;
#10000;
data_in <= 24'b000010000000101100001001;
#10000;
data_in <= 24'b010100010110011010000010;
#10000;
data_in <= 24'b001111110101001001100111;
#10000;
data_in <= 24'b000110000010011100110111;
#10000;
data_in <= 24'b000000010000101100010101;
#10000;
data_in <= 24'b000010000000111000010011;
#10000;
data_in <= 24'b000010010000111000001111;
#10000;
data_in <= 24'b000001010000100000000110;
#10000;
data_in <= 24'b000010100000101100000111;
#10000;
data_in <= 24'b010100000110010110000000;
#10000;
data_in <= 24'b010000000101001101101000;
#10000;
data_in <= 24'b000110100010011100110111;
#10000;
data_in <= 24'b000000000000100100010001;
#10000;
data_in <= 24'b000000110000101000001101;
#10000;
data_in <= 24'b000001000000100100001000;
#10000;
data_in <= 24'b000001000000011100000101;
#10000;
data_in <= 24'b000100010001001000001110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000111000010011000111000;
#10000;
data_in <= 24'b000100010001101100101101;
#10000;
data_in <= 24'b000011000001011000100111;
#10000;
data_in <= 24'b000101000001111000101111;
#10000;
data_in <= 24'b000111010010011000110100;
#10000;
data_in <= 24'b000111000010010100110011;
#10000;
data_in <= 24'b000110000010000100101111;
#10000;
data_in <= 24'b000101010001111100110000;
#10000;
data_in <= 24'b000101000001111000110000;
#10000;
data_in <= 24'b000011000001011000101000;
#10000;
data_in <= 24'b000010100001010000100101;
#10000;
data_in <= 24'b000101000001111000101111;
#10000;
data_in <= 24'b000111100010011100110101;
#10000;
data_in <= 24'b000111010010011000110100;
#10000;
data_in <= 24'b000110110010010000110010;
#10000;
data_in <= 24'b000110110010010000110010;
#10000;
data_in <= 24'b000011010001011100101001;
#10000;
data_in <= 24'b000010000001001000100100;
#10000;
data_in <= 24'b000011010001010100100110;
#10000;
data_in <= 24'b000101110001111100110000;
#10000;
data_in <= 24'b000111100010010100110100;
#10000;
data_in <= 24'b000111000010010000110001;
#10000;
data_in <= 24'b000110110010001100110000;
#10000;
data_in <= 24'b000111010010011000110011;
#10000;
data_in <= 24'b000011000001011000101000;
#10000;
data_in <= 24'b000010010001001100100101;
#10000;
data_in <= 24'b000011110001011100101000;
#10000;
data_in <= 24'b000110000010000100101111;
#10000;
data_in <= 24'b000111000010001100110010;
#10000;
data_in <= 24'b000110000010000000101101;
#10000;
data_in <= 24'b000101110001111100101100;
#10000;
data_in <= 24'b000111000010010000110001;
#10000;
data_in <= 24'b000011000001010100101001;
#10000;
data_in <= 24'b000010010001001100100101;
#10000;
data_in <= 24'b000011100001011000100111;
#10000;
data_in <= 24'b000101100001111100101101;
#10000;
data_in <= 24'b000110000001111100101110;
#10000;
data_in <= 24'b000101100001110000101001;
#10000;
data_in <= 24'b000101100001110000100111;
#10000;
data_in <= 24'b000111000010001000101101;
#10000;
data_in <= 24'b000011110001100000101100;
#10000;
data_in <= 24'b000010100001010000100110;
#10000;
data_in <= 24'b000011000001001100100110;
#10000;
data_in <= 24'b000100100001100100101000;
#10000;
data_in <= 24'b000101100001110000101001;
#10000;
data_in <= 24'b000100110001100100100100;
#10000;
data_in <= 24'b000101110001110000100101;
#10000;
data_in <= 24'b000111010010001000101011;
#10000;
data_in <= 24'b000101110010000000110100;
#10000;
data_in <= 24'b000011100001100000101010;
#10000;
data_in <= 24'b000010110001001000100101;
#10000;
data_in <= 24'b000011110001011000100101;
#10000;
data_in <= 24'b000100100001100000100101;
#10000;
data_in <= 24'b000100010001010100100000;
#10000;
data_in <= 24'b000101010001011100100001;
#10000;
data_in <= 24'b000110000001110100100110;
#10000;
data_in <= 24'b001000010010100000111011;
#10000;
data_in <= 24'b000101010001110000101111;
#10000;
data_in <= 24'b000011000001010000100101;
#10000;
data_in <= 24'b000011010001010000100011;
#10000;
data_in <= 24'b000011100001010000011111;
#10000;
data_in <= 24'b000011010001001000011011;
#10000;
data_in <= 24'b000011010001001000011011;
#10000;
data_in <= 24'b000100000001011100100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000010100001011100100111;
#10000;
data_in <= 24'b000000000000110000011110;
#10000;
data_in <= 24'b000011010001101100110001;
#10000;
data_in <= 24'b001110010100100101100000;
#10000;
data_in <= 24'b010100010110010001111111;
#10000;
data_in <= 24'b010010010101111001111001;
#10000;
data_in <= 24'b001111000101001001101110;
#10000;
data_in <= 24'b001111010101001001101110;
#10000;
data_in <= 24'b000011110001100100101010;
#10000;
data_in <= 24'b000000100000111100011111;
#10000;
data_in <= 24'b000010000001011000101001;
#10000;
data_in <= 24'b001010010011101001001111;
#10000;
data_in <= 24'b010001110101100001110010;
#10000;
data_in <= 24'b010010110101111001111001;
#10000;
data_in <= 24'b010000100101011101110010;
#10000;
data_in <= 24'b001111010101010001101110;
#10000;
data_in <= 24'b000101000001110100101011;
#10000;
data_in <= 24'b000001110001000100100010;
#10000;
data_in <= 24'b000000100001000000100010;
#10000;
data_in <= 24'b000101100010010100111000;
#10000;
data_in <= 24'b001101010100010101011100;
#10000;
data_in <= 24'b010001110101101101110100;
#10000;
data_in <= 24'b010001110101110001110111;
#10000;
data_in <= 24'b001111110101011001110000;
#10000;
data_in <= 24'b000101010001110100101010;
#10000;
data_in <= 24'b000011000001011100100101;
#10000;
data_in <= 24'b000000110001000000100000;
#10000;
data_in <= 24'b000001110001011100101000;
#10000;
data_in <= 24'b001000010011001001000111;
#10000;
data_in <= 24'b001111010101001001101000;
#10000;
data_in <= 24'b010010000101111001110111;
#10000;
data_in <= 24'b010001000101101101110101;
#10000;
data_in <= 24'b000100110001110000100110;
#10000;
data_in <= 24'b000100010001101000100111;
#10000;
data_in <= 24'b000010100001010000100101;
#10000;
data_in <= 24'b000001010001001100100101;
#10000;
data_in <= 24'b000101000010010100111010;
#10000;
data_in <= 24'b001011010100001001011000;
#10000;
data_in <= 24'b010000010101011101110000;
#10000;
data_in <= 24'b010001110101111001111000;
#10000;
data_in <= 24'b000100110001100100100100;
#10000;
data_in <= 24'b000100000001101000100100;
#10000;
data_in <= 24'b000011100001100100100111;
#10000;
data_in <= 24'b000010110001100100101011;
#10000;
data_in <= 24'b000011110010000000110011;
#10000;
data_in <= 24'b000111000011000101000111;
#10000;
data_in <= 24'b001100100100100001100001;
#10000;
data_in <= 24'b010000110101101001110100;
#10000;
data_in <= 24'b000100100001100100100010;
#10000;
data_in <= 24'b000011000001010100011111;
#10000;
data_in <= 24'b000011100001100100100111;
#10000;
data_in <= 24'b000100110010001000110010;
#10000;
data_in <= 24'b000100010010001000110101;
#10000;
data_in <= 24'b000011110010010000111010;
#10000;
data_in <= 24'b001000000011011001001111;
#10000;
data_in <= 24'b001110010101000001101010;
#10000;
data_in <= 24'b000100000001100100100010;
#10000;
data_in <= 24'b000001110001001000011010;
#10000;
data_in <= 24'b000011000001100000100100;
#10000;
data_in <= 24'b000110010010100100110110;
#10000;
data_in <= 24'b000101010010011100111000;
#10000;
data_in <= 24'b000010100001110100110010;
#10000;
data_in <= 24'b000101110010110001000010;
#10000;
data_in <= 24'b001100010100011101100000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001111000101000001101001;
#10000;
data_in <= 24'b010000110101010001101110;
#10000;
data_in <= 24'b010000110101010001101110;
#10000;
data_in <= 24'b010001000101010101101111;
#10000;
data_in <= 24'b010001010101011001110000;
#10000;
data_in <= 24'b001111000100110101100111;
#10000;
data_in <= 24'b001101110100100001100011;
#10000;
data_in <= 24'b001110110100111001101001;
#10000;
data_in <= 24'b010000100101011101110010;
#10000;
data_in <= 24'b010010010101110001110111;
#10000;
data_in <= 24'b010010010101110001110111;
#10000;
data_in <= 24'b010010100101110001111001;
#10000;
data_in <= 24'b010011000101111001111011;
#10000;
data_in <= 24'b010001000101100101110101;
#10000;
data_in <= 24'b010000100101011001110101;
#10000;
data_in <= 24'b010010100101111001111101;
#10000;
data_in <= 24'b010010000101110101111000;
#10000;
data_in <= 24'b010011000110000101111101;
#10000;
data_in <= 24'b010010110110000001111100;
#10000;
data_in <= 24'b010011010110000110000000;
#10000;
data_in <= 24'b010100100110011010000101;
#10000;
data_in <= 24'b010011100110001110000011;
#10000;
data_in <= 24'b010011110110001110000110;
#10000;
data_in <= 24'b010110000110111010010001;
#10000;
data_in <= 24'b010010000101110101111001;
#10000;
data_in <= 24'b010011000110000101111101;
#10000;
data_in <= 24'b010010110101111101111110;
#10000;
data_in <= 24'b010011000110000110000001;
#10000;
data_in <= 24'b010100100110011110000111;
#10000;
data_in <= 24'b010100000110011010001001;
#10000;
data_in <= 24'b010101000110101010001110;
#10000;
data_in <= 24'b010111100111010110011011;
#10000;
data_in <= 24'b010010000101111001111010;
#10000;
data_in <= 24'b010010110110000001111111;
#10000;
data_in <= 24'b010010100101111101111111;
#10000;
data_in <= 24'b010010100110000110000001;
#10000;
data_in <= 24'b010100010110011110001011;
#10000;
data_in <= 24'b010100000110011110001101;
#10000;
data_in <= 24'b010100100110101110010011;
#10000;
data_in <= 24'b010111100111100010100000;
#10000;
data_in <= 24'b010010000101110101111100;
#10000;
data_in <= 24'b010010100110001010000000;
#10000;
data_in <= 24'b010010100110000110000001;
#10000;
data_in <= 24'b010010110110010010000110;
#10000;
data_in <= 24'b010100100110100110001111;
#10000;
data_in <= 24'b010100010110101010010010;
#10000;
data_in <= 24'b010101000110110110010111;
#10000;
data_in <= 24'b010111100111101010100011;
#10000;
data_in <= 24'b010000010101100101110111;
#10000;
data_in <= 24'b010001110101111101111101;
#10000;
data_in <= 24'b010010010110000010000000;
#10000;
data_in <= 24'b010011000110010110000111;
#10000;
data_in <= 24'b010101000110101110010001;
#10000;
data_in <= 24'b010100100110101110010011;
#10000;
data_in <= 24'b010101000110110110010111;
#10000;
data_in <= 24'b010111010111100010100100;
#10000;
data_in <= 24'b001111010101001101101111;
#10000;
data_in <= 24'b010000100101101001111000;
#10000;
data_in <= 24'b010001010101110001111100;
#10000;
data_in <= 24'b010010010110001010000100;
#10000;
data_in <= 24'b010100100110100110001111;
#10000;
data_in <= 24'b010100000110100110010001;
#10000;
data_in <= 24'b010100010110101010010100;
#10000;
data_in <= 24'b010110110111011010100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010010110110000001111100;
#10000;
data_in <= 24'b011001000111100110011000;
#10000;
data_in <= 24'b100001101001110110111101;
#10000;
data_in <= 24'b101000101011101111011101;
#10000;
data_in <= 24'b101101001100111111110001;
#10000;
data_in <= 24'b101110111101011111111010;
#10000;
data_in <= 24'b101110001101001111111000;
#10000;
data_in <= 24'b101011101100111011110001;
#10000;
data_in <= 24'b011000100111011110010111;
#10000;
data_in <= 24'b011110001000111110101111;
#10000;
data_in <= 24'b100101001010110111001111;
#10000;
data_in <= 24'b101010011100001111100111;
#10000;
data_in <= 24'b101101011101000111110100;
#10000;
data_in <= 24'b101110001101011011111001;
#10000;
data_in <= 24'b101101111101010011111001;
#10000;
data_in <= 24'b101100011101000111110101;
#10000;
data_in <= 24'b011101001000110010110000;
#10000;
data_in <= 24'b100001111010000111000101;
#10000;
data_in <= 24'b101000001011101011011110;
#10000;
data_in <= 24'b101011101100100111101110;
#10000;
data_in <= 24'b101100101100111111110100;
#10000;
data_in <= 24'b101101001101010011111000;
#10000;
data_in <= 24'b101101011101010111111001;
#10000;
data_in <= 24'b101100101101010011111000;
#10000;
data_in <= 24'b011101101000111110110111;
#10000;
data_in <= 24'b100010101010010011001100;
#10000;
data_in <= 24'b101000011011101111100011;
#10000;
data_in <= 24'b101010111100100011101101;
#10000;
data_in <= 24'b101011011100110111110001;
#10000;
data_in <= 24'b101100001101000011110100;
#10000;
data_in <= 24'b101100111101001111110111;
#10000;
data_in <= 24'b101100111101010111111001;
#10000;
data_in <= 24'b011101011000111010111000;
#10000;
data_in <= 24'b100001111010001111001100;
#10000;
data_in <= 24'b100111111011101111100100;
#10000;
data_in <= 24'b101010011100100011101111;
#10000;
data_in <= 24'b101011011100110011110011;
#10000;
data_in <= 24'b101011011100111011110101;
#10000;
data_in <= 24'b101011111101000111110101;
#10000;
data_in <= 24'b101100001101001011110110;
#10000;
data_in <= 24'b011101101001000110111101;
#10000;
data_in <= 24'b100010001010010111010001;
#10000;
data_in <= 24'b100111101011101111100111;
#10000;
data_in <= 24'b101010001100100011110001;
#10000;
data_in <= 24'b101011001100110111110100;
#10000;
data_in <= 24'b101011101100111111110110;
#10000;
data_in <= 24'b101011011100111111110011;
#10000;
data_in <= 24'b101011001100111011110010;
#10000;
data_in <= 24'b011101111001000110111111;
#10000;
data_in <= 24'b100001101010001111001111;
#10000;
data_in <= 24'b100110101011011111100011;
#10000;
data_in <= 24'b101001011100010111101110;
#10000;
data_in <= 24'b101010101100101111110010;
#10000;
data_in <= 24'b101010101100111011110100;
#10000;
data_in <= 24'b101010001100110011110000;
#10000;
data_in <= 24'b101001011100100111101101;
#10000;
data_in <= 24'b011100101000111110111011;
#10000;
data_in <= 24'b100000101001111111001100;
#10000;
data_in <= 24'b100100101011001011011101;
#10000;
data_in <= 24'b100111001011111011101001;
#10000;
data_in <= 24'b101001001100011111101111;
#10000;
data_in <= 24'b101001101100101111110001;
#10000;
data_in <= 24'b101001011100101011110000;
#10000;
data_in <= 24'b101000101100011011101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101011011101001111110011;
#10000;
data_in <= 24'b101011001101010111110101;
#10000;
data_in <= 24'b101010111101010011110100;
#10000;
data_in <= 24'b101010001101000111110010;
#10000;
data_in <= 24'b101001111100111111110010;
#10000;
data_in <= 24'b101000111100101111101110;
#10000;
data_in <= 24'b100110111011111111100111;
#10000;
data_in <= 24'b100011111011001111011011;
#10000;
data_in <= 24'b101011101101010011110110;
#10000;
data_in <= 24'b101011011101011011110110;
#10000;
data_in <= 24'b101011001101010111110110;
#10000;
data_in <= 24'b101010011101001011110011;
#10000;
data_in <= 24'b101010001101000011110011;
#10000;
data_in <= 24'b101001001100110011101111;
#10000;
data_in <= 24'b100111001100000111100111;
#10000;
data_in <= 24'b100100011011010111011101;
#10000;
data_in <= 24'b101100001101010111110111;
#10000;
data_in <= 24'b101100001101011011111000;
#10000;
data_in <= 24'b101011111101010111110111;
#10000;
data_in <= 24'b101011011101001111110101;
#10000;
data_in <= 24'b101010111101000111110100;
#10000;
data_in <= 24'b101001111100110111110000;
#10000;
data_in <= 24'b101000001100010011101010;
#10000;
data_in <= 24'b100101111011101111100001;
#10000;
data_in <= 24'b101100011101011011111000;
#10000;
data_in <= 24'b101100001101011011111000;
#10000;
data_in <= 24'b101011111101010111110111;
#10000;
data_in <= 24'b101011101101010011110110;
#10000;
data_in <= 24'b101011001101001011110101;
#10000;
data_in <= 24'b101010001100111011110001;
#10000;
data_in <= 24'b101000101100011011101100;
#10000;
data_in <= 24'b100111011100000111100111;
#10000;
data_in <= 24'b101011111101001111110111;
#10000;
data_in <= 24'b101011111101001111110111;
#10000;
data_in <= 24'b101011111101001111110111;
#10000;
data_in <= 24'b101011111101001111110111;
#10000;
data_in <= 24'b101011011101000111110101;
#10000;
data_in <= 24'b101010011100110111110001;
#10000;
data_in <= 24'b101001111100100011101111;
#10000;
data_in <= 24'b101001001100010111101100;
#10000;
data_in <= 24'b101011001101000011110100;
#10000;
data_in <= 24'b101010111100111111110011;
#10000;
data_in <= 24'b101011001101000011110100;
#10000;
data_in <= 24'b101011101101001011110110;
#10000;
data_in <= 24'b101011001101000011110100;
#10000;
data_in <= 24'b101010011100110111110001;
#10000;
data_in <= 24'b101010001100100111110000;
#10000;
data_in <= 24'b101010011100101011110001;
#10000;
data_in <= 24'b101010111100110111110001;
#10000;
data_in <= 24'b101010011100101111101111;
#10000;
data_in <= 24'b101010101100110011110000;
#10000;
data_in <= 24'b101011101101000011110100;
#10000;
data_in <= 24'b101011011100111111110011;
#10000;
data_in <= 24'b101010011100101111101111;
#10000;
data_in <= 24'b101010011100101011110001;
#10000;
data_in <= 24'b101011001100110111110100;
#10000;
data_in <= 24'b101001101100101011110000;
#10000;
data_in <= 24'b101001001100100011101110;
#10000;
data_in <= 24'b101010001100100111110000;
#10000;
data_in <= 24'b101010101100111011110010;
#10000;
data_in <= 24'b101011001100111011110010;
#10000;
data_in <= 24'b101001111100101111101111;
#10000;
data_in <= 24'b101010001100110011110000;
#10000;
data_in <= 24'b101011001101000011110100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100010001010101011010101;
#10000;
data_in <= 24'b011111111010000111001100;
#10000;
data_in <= 24'b011011101000111010111001;
#10000;
data_in <= 24'b010010000110010110010001;
#10000;
data_in <= 24'b000011110010101001010110;
#10000;
data_in <= 24'b000000000000010100101111;
#10000;
data_in <= 24'b000000000001010000111110;
#10000;
data_in <= 24'b001000000011100101100011;
#10000;
data_in <= 24'b100000111010010111010000;
#10000;
data_in <= 24'b011110011001101111000110;
#10000;
data_in <= 24'b011001001000010010101111;
#10000;
data_in <= 24'b001111100101101110000111;
#10000;
data_in <= 24'b000100010010110001011000;
#10000;
data_in <= 24'b000000000001001100111111;
#10000;
data_in <= 24'b000010010010001001001110;
#10000;
data_in <= 24'b001001100011111101101001;
#10000;
data_in <= 24'b100000001010001111001011;
#10000;
data_in <= 24'b011001111000101010110010;
#10000;
data_in <= 24'b010011100110111010011001;
#10000;
data_in <= 24'b001101100101001101111111;
#10000;
data_in <= 24'b000101100011001101011111;
#10000;
data_in <= 24'b000001010010000001001100;
#10000;
data_in <= 24'b000101100011000101011101;
#10000;
data_in <= 24'b001110000101001101111111;
#10000;
data_in <= 24'b100100101011010111011101;
#10000;
data_in <= 24'b011010001000101110110011;
#10000;
data_in <= 24'b010010010110100110010100;
#10000;
data_in <= 24'b001111010101110110001000;
#10000;
data_in <= 24'b001010100100101001110101;
#10000;
data_in <= 24'b000111010011101001100110;
#10000;
data_in <= 24'b001110010101011010000011;
#10000;
data_in <= 24'b011010011000011010110011;
#10000;
data_in <= 24'b100111001011110011100101;
#10000;
data_in <= 24'b011110001001100011000001;
#10000;
data_in <= 24'b010011110110111110011010;
#10000;
data_in <= 24'b001101100101011010000001;
#10000;
data_in <= 24'b001010100100100101110110;
#10000;
data_in <= 24'b001101100101010110000010;
#10000;
data_in <= 24'b011000000111111010101101;
#10000;
data_in <= 24'b100011001010101011011001;
#10000;
data_in <= 24'b100111011011110111100110;
#10000;
data_in <= 24'b100100001011000011011001;
#10000;
data_in <= 24'b011010011000100110110100;
#10000;
data_in <= 24'b001110100101110010000111;
#10000;
data_in <= 24'b001101000101010110000010;
#10000;
data_in <= 24'b010110010111101010100111;
#10000;
data_in <= 24'b100000111010010011010010;
#10000;
data_in <= 24'b100101101011011111100101;
#10000;
data_in <= 24'b101010111100101111110100;
#10000;
data_in <= 24'b101010111100101111110100;
#10000;
data_in <= 24'b100101001011011011100001;
#10000;
data_in <= 24'b011101101001100011000011;
#10000;
data_in <= 24'b011100111001010011000001;
#10000;
data_in <= 24'b100010111010111011011010;
#10000;
data_in <= 24'b100111011011111111101101;
#10000;
data_in <= 24'b100111001011110111101011;
#10000;
data_in <= 24'b101010011100110111110011;
#10000;
data_in <= 24'b101001011100100011110000;
#10000;
data_in <= 24'b101001001100011111101111;
#10000;
data_in <= 24'b101001101100100111110100;
#10000;
data_in <= 24'b101001101100100111110101;
#10000;
data_in <= 24'b100111011100000111101111;
#10000;
data_in <= 24'b100101011011011011100111;
#10000;
data_in <= 24'b100011111011000011100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101100101001001111011;
#10000;
data_in <= 24'b001010110100100101110010;
#10000;
data_in <= 24'b001001110100010001110000;
#10000;
data_in <= 24'b001111000101100110000101;
#10000;
data_in <= 24'b011010011000100010110101;
#10000;
data_in <= 24'b100100111011010011100010;
#10000;
data_in <= 24'b100111111011111111110000;
#10000;
data_in <= 24'b100101101011011111101000;
#10000;
data_in <= 24'b001011010100100101110010;
#10000;
data_in <= 24'b001101110101010010000000;
#10000;
data_in <= 24'b010010110110100010010100;
#10000;
data_in <= 24'b011010111000100010110101;
#10000;
data_in <= 24'b100100001010111011011101;
#10000;
data_in <= 24'b101010111100100111111010;
#10000;
data_in <= 24'b101001111100011011111001;
#10000;
data_in <= 24'b100101111011011111101100;
#10000;
data_in <= 24'b010110010111011010100010;
#10000;
data_in <= 24'b011010001000010110110001;
#10000;
data_in <= 24'b011110111001100011000101;
#10000;
data_in <= 24'b100011111010101111011010;
#10000;
data_in <= 24'b101000001011111011101111;
#10000;
data_in <= 24'b101011011100101011111101;
#10000;
data_in <= 24'b101001111100011011111011;
#10000;
data_in <= 24'b100110111011101011110001;
#10000;
data_in <= 24'b100101101011001111100000;
#10000;
data_in <= 24'b100111001011100111100110;
#10000;
data_in <= 24'b100111111011101111101010;
#10000;
data_in <= 24'b100111111011101011101100;
#10000;
data_in <= 24'b100111101011101111101110;
#10000;
data_in <= 24'b101000001011110011110010;
#10000;
data_in <= 24'b100111001011101011110001;
#10000;
data_in <= 24'b100101111011010011101101;
#10000;
data_in <= 24'b101001011100001111110010;
#10000;
data_in <= 24'b101010001100011011110101;
#10000;
data_in <= 24'b101010111100100111111000;
#10000;
data_in <= 24'b101010011100011111111000;
#10000;
data_in <= 24'b101001011100000111110111;
#10000;
data_in <= 24'b100111001011011111101111;
#10000;
data_in <= 24'b100100001010101011100110;
#10000;
data_in <= 24'b100001101010000011011100;
#10000;
data_in <= 24'b101000111100000111110000;
#10000;
data_in <= 24'b101000111100000111110010;
#10000;
data_in <= 24'b101000111100000111110010;
#10000;
data_in <= 24'b101000101011111111110010;
#10000;
data_in <= 24'b100111011011100011110000;
#10000;
data_in <= 24'b100100011010110011100101;
#10000;
data_in <= 24'b100000001001100111010111;
#10000;
data_in <= 24'b011100111000110011001100;
#10000;
data_in <= 24'b100111101011110011101101;
#10000;
data_in <= 24'b100110001011011011100111;
#10000;
data_in <= 24'b100011111010110011011111;
#10000;
data_in <= 24'b100010001010010011011010;
#10000;
data_in <= 24'b100000101001110111010101;
#10000;
data_in <= 24'b011110101001010111001110;
#10000;
data_in <= 24'b011100101000100111000111;
#10000;
data_in <= 24'b011011001000001011000011;
#10000;
data_in <= 24'b100011101010110011100011;
#10000;
data_in <= 24'b100010001010001111011100;
#10000;
data_in <= 24'b011111101001100011010100;
#10000;
data_in <= 24'b011101111001000011001110;
#10000;
data_in <= 24'b011100101000100111000111;
#10000;
data_in <= 24'b011011011000001111000100;
#10000;
data_in <= 24'b011010110111111011000001;
#10000;
data_in <= 24'b011010010111110010111111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100101001011011111101001;
#10000;
data_in <= 24'b100101001011100011101000;
#10000;
data_in <= 24'b100100101011100011101000;
#10000;
data_in <= 24'b100100101011100011101000;
#10000;
data_in <= 24'b100100101011101011101010;
#10000;
data_in <= 24'b100101001011110111101010;
#10000;
data_in <= 24'b100101011011111111101100;
#10000;
data_in <= 24'b100101101100000011101101;
#10000;
data_in <= 24'b100101111011011111101100;
#10000;
data_in <= 24'b100101001011011011101011;
#10000;
data_in <= 24'b100100011011001111101000;
#10000;
data_in <= 24'b100011011011001011100110;
#10000;
data_in <= 24'b100011011011001011100100;
#10000;
data_in <= 24'b100011011011010111100110;
#10000;
data_in <= 24'b100011111011011111101000;
#10000;
data_in <= 24'b100100011011100111101010;
#10000;
data_in <= 24'b100100101011000111101000;
#10000;
data_in <= 24'b100011011010111111100101;
#10000;
data_in <= 24'b100010011010101011100010;
#10000;
data_in <= 24'b100001011010011011011110;
#10000;
data_in <= 24'b100001001010011011011100;
#10000;
data_in <= 24'b100000111010011111011101;
#10000;
data_in <= 24'b100001011010100111011111;
#10000;
data_in <= 24'b100010011010101111100001;
#10000;
data_in <= 24'b100000101001111011011010;
#10000;
data_in <= 24'b011111101001110011010111;
#10000;
data_in <= 24'b011110101001011111010100;
#10000;
data_in <= 24'b011101101001001111010000;
#10000;
data_in <= 24'b011101001001001011001101;
#10000;
data_in <= 24'b011100111001000111001100;
#10000;
data_in <= 24'b011101001001001011001101;
#10000;
data_in <= 24'b011101011001001111001110;
#10000;
data_in <= 24'b011101101000111111001101;
#10000;
data_in <= 24'b011100101000111011001011;
#10000;
data_in <= 24'b011011011000100011001000;
#10000;
data_in <= 24'b011010001000001111000011;
#10000;
data_in <= 24'b011000110111111010111110;
#10000;
data_in <= 24'b010111110111101010111010;
#10000;
data_in <= 24'b010111000111011110110111;
#10000;
data_in <= 24'b010110110111011010110110;
#10000;
data_in <= 24'b011101011000111011001110;
#10000;
data_in <= 24'b011100011000100111001011;
#10000;
data_in <= 24'b011010111000001111000101;
#10000;
data_in <= 24'b011000100111101010111100;
#10000;
data_in <= 24'b010111000111000110110101;
#10000;
data_in <= 24'b010101000110110010101110;
#10000;
data_in <= 24'b010100010110011010101010;
#10000;
data_in <= 24'b010011010110010110100111;
#10000;
data_in <= 24'b011100001000011011001000;
#10000;
data_in <= 24'b011010100111111111000011;
#10000;
data_in <= 24'b011000010111011010111010;
#10000;
data_in <= 24'b010101100110101110101111;
#10000;
data_in <= 24'b010100000110001010101001;
#10000;
data_in <= 24'b010010000101110110100001;
#10000;
data_in <= 24'b010010000101101010100001;
#10000;
data_in <= 24'b010001100101101110011111;
#10000;
data_in <= 24'b011000100111010110111001;
#10000;
data_in <= 24'b010111000110110010110001;
#10000;
data_in <= 24'b010100010110000110100110;
#10000;
data_in <= 24'b010001100101011010011011;
#10000;
data_in <= 24'b001111110101000010010011;
#10000;
data_in <= 24'b001111010100111010010001;
#10000;
data_in <= 24'b001111110101000010010011;
#10000;
data_in <= 24'b010000000101000110010100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100101001011101111101000;
#10000;
data_in <= 24'b100100111011101011100111;
#10000;
data_in <= 24'b100100111011011111100101;
#10000;
data_in <= 24'b100100011011010111100011;
#10000;
data_in <= 24'b100011111011001111100001;
#10000;
data_in <= 24'b100010111010111111011101;
#10000;
data_in <= 24'b100010011010110011011000;
#10000;
data_in <= 24'b100001101010100111010101;
#10000;
data_in <= 24'b100100001011010111100111;
#10000;
data_in <= 24'b100100101011010111100111;
#10000;
data_in <= 24'b100100001011001111100101;
#10000;
data_in <= 24'b100011111011001111100011;
#10000;
data_in <= 24'b100011011011000111100001;
#10000;
data_in <= 24'b100010011010110111011011;
#10000;
data_in <= 24'b100001111010100111010111;
#10000;
data_in <= 24'b100001001010011111010011;
#10000;
data_in <= 24'b100010001010101011100000;
#10000;
data_in <= 24'b100011001010101111100010;
#10000;
data_in <= 24'b100011101010111011100011;
#10000;
data_in <= 24'b100011111010111111100100;
#10000;
data_in <= 24'b100011101010111111100001;
#10000;
data_in <= 24'b100010101010101111011100;
#10000;
data_in <= 24'b100001101010100011010110;
#10000;
data_in <= 24'b100000111010011011010010;
#10000;
data_in <= 24'b011101101001010011001111;
#10000;
data_in <= 24'b011111001001101011010011;
#10000;
data_in <= 24'b100000111010000111011010;
#10000;
data_in <= 24'b100010011010100011011111;
#10000;
data_in <= 24'b100010101010101011011111;
#10000;
data_in <= 24'b100010001010100111011011;
#10000;
data_in <= 24'b100001001010010111010110;
#10000;
data_in <= 24'b100000011010001111010001;
#10000;
data_in <= 24'b010111000111100010110101;
#10000;
data_in <= 24'b011000110111111110111100;
#10000;
data_in <= 24'b011011101000101011000111;
#10000;
data_in <= 24'b011101101001001011001110;
#10000;
data_in <= 24'b011110111001100111010000;
#10000;
data_in <= 24'b011111011001110011010001;
#10000;
data_in <= 24'b011111101001111011001111;
#10000;
data_in <= 24'b011111111010000011001110;
#10000;
data_in <= 24'b010001110101111110100001;
#10000;
data_in <= 24'b010010010110010010100100;
#10000;
data_in <= 24'b010011100110100110101001;
#10000;
data_in <= 24'b010101000111000010101100;
#10000;
data_in <= 24'b010110110111100010110001;
#10000;
data_in <= 24'b011001111000011010111011;
#10000;
data_in <= 24'b011101001001001111000110;
#10000;
data_in <= 24'b011111011001110111001110;
#10000;
data_in <= 24'b010000000101010110011001;
#10000;
data_in <= 24'b001110010101000110010011;
#10000;
data_in <= 24'b001100100100101110001011;
#10000;
data_in <= 24'b001100000100100110000111;
#10000;
data_in <= 24'b001110100101010010010000;
#10000;
data_in <= 24'b010100010110110010100100;
#10000;
data_in <= 24'b011011001000101111000000;
#10000;
data_in <= 24'b100000011010000111010010;
#10000;
data_in <= 24'b010000110101010110011100;
#10000;
data_in <= 24'b001101000100100110001101;
#10000;
data_in <= 24'b001000110011100101111011;
#10000;
data_in <= 24'b000110100011000001110001;
#10000;
data_in <= 24'b001000100011110001111000;
#10000;
data_in <= 24'b010000100101110110010110;
#10000;
data_in <= 24'b011010011000100010111101;
#10000;
data_in <= 24'b100001101010011011010111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100000001010001011001101;
#10000;
data_in <= 24'b011111001001111011001001;
#10000;
data_in <= 24'b011110011001100111000100;
#10000;
data_in <= 24'b011101011001010111000000;
#10000;
data_in <= 24'b011100101001001010111011;
#10000;
data_in <= 24'b011011111000111110111000;
#10000;
data_in <= 24'b011011111000110110110110;
#10000;
data_in <= 24'b011011001000110010110111;
#10000;
data_in <= 24'b100000101010010011001111;
#10000;
data_in <= 24'b011111101010000011001011;
#10000;
data_in <= 24'b011110111001101111000110;
#10000;
data_in <= 24'b011101101001011011000001;
#10000;
data_in <= 24'b011100101001001010111011;
#10000;
data_in <= 24'b011011111000111110111000;
#10000;
data_in <= 24'b011010111000101110110100;
#10000;
data_in <= 24'b011001111000100010110101;
#10000;
data_in <= 24'b100000111010010111010000;
#10000;
data_in <= 24'b100000001010001011001101;
#10000;
data_in <= 24'b011110111001110111001000;
#10000;
data_in <= 24'b011101101001100011000011;
#10000;
data_in <= 24'b011100011001001110111110;
#10000;
data_in <= 24'b011011001000111010111001;
#10000;
data_in <= 24'b011001111000100110110100;
#10000;
data_in <= 24'b011000111000011010110010;
#10000;
data_in <= 24'b100000101010001111010000;
#10000;
data_in <= 24'b011111111010000111001100;
#10000;
data_in <= 24'b011110111001110111001000;
#10000;
data_in <= 24'b011101101001100011000011;
#10000;
data_in <= 24'b011100101001010010111111;
#10000;
data_in <= 24'b011011011000111110111010;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011000111000011010110010;
#10000;
data_in <= 24'b011111101010000111001101;
#10000;
data_in <= 24'b011110111001111011001010;
#10000;
data_in <= 24'b011110001001101111000111;
#10000;
data_in <= 24'b011101001001011111000011;
#10000;
data_in <= 24'b011100011001010011000000;
#10000;
data_in <= 24'b011011011001000010111100;
#10000;
data_in <= 24'b011010001000101110110111;
#10000;
data_in <= 24'b011000111000100010110100;
#10000;
data_in <= 24'b011111001001111011001100;
#10000;
data_in <= 24'b011110011001110011001000;
#10000;
data_in <= 24'b011101011001100011000100;
#10000;
data_in <= 24'b011100101001010111000001;
#10000;
data_in <= 24'b011011111001001010111110;
#10000;
data_in <= 24'b011011001000111110111011;
#10000;
data_in <= 24'b011010011000110010111000;
#10000;
data_in <= 24'b011001001000100110110101;
#10000;
data_in <= 24'b011110111001110111001011;
#10000;
data_in <= 24'b011110001001101011001000;
#10000;
data_in <= 24'b011100011001011011000010;
#10000;
data_in <= 24'b011011101001001110111111;
#10000;
data_in <= 24'b011010111000111110111101;
#10000;
data_in <= 24'b011010001000110010111010;
#10000;
data_in <= 24'b011001101000101010111000;
#10000;
data_in <= 24'b011000101000100110110101;
#10000;
data_in <= 24'b011111001001111011001100;
#10000;
data_in <= 24'b011110001001101111000111;
#10000;
data_in <= 24'b011100011001011011000010;
#10000;
data_in <= 24'b011011001001001010111100;
#10000;
data_in <= 24'b011010011000111010111010;
#10000;
data_in <= 24'b011001111000110010111000;
#10000;
data_in <= 24'b011001001000100110110101;
#10000;
data_in <= 24'b011000011000100110110011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011001001000011110111001;
#10000;
data_in <= 24'b011000001000010110111001;
#10000;
data_in <= 24'b010111111000001010110100;
#10000;
data_in <= 24'b010111111000000110101111;
#10000;
data_in <= 24'b010111100111111110101100;
#10000;
data_in <= 24'b010111010111101110100100;
#10000;
data_in <= 24'b010110100111010110011010;
#10000;
data_in <= 24'b010110000111000110010001;
#10000;
data_in <= 24'b011001101000101010111010;
#10000;
data_in <= 24'b011000101000011110111001;
#10000;
data_in <= 24'b011000011000010110110101;
#10000;
data_in <= 24'b011000011000001110110001;
#10000;
data_in <= 24'b011000001000000110101110;
#10000;
data_in <= 24'b010111110111110110100110;
#10000;
data_in <= 24'b010111000111100010011011;
#10000;
data_in <= 24'b010110010111001110010001;
#10000;
data_in <= 24'b011001011000101110111011;
#10000;
data_in <= 24'b011000101000100010111000;
#10000;
data_in <= 24'b011000101000011010110110;
#10000;
data_in <= 24'b011000101000010110110001;
#10000;
data_in <= 24'b011000001000001010101101;
#10000;
data_in <= 24'b010111010111111010100101;
#10000;
data_in <= 24'b010110110111011110011010;
#10000;
data_in <= 24'b010110000111001010010000;
#10000;
data_in <= 24'b011000111000101010110111;
#10000;
data_in <= 24'b010111111000100010110101;
#10000;
data_in <= 24'b010111101000010110110010;
#10000;
data_in <= 24'b010111101000001110101111;
#10000;
data_in <= 24'b010111101000001010101010;
#10000;
data_in <= 24'b010110100111101110100010;
#10000;
data_in <= 24'b010110000111010010010111;
#10000;
data_in <= 24'b010101010110111110001101;
#10000;
data_in <= 24'b011000101000100110110101;
#10000;
data_in <= 24'b010111101000100010110011;
#10000;
data_in <= 24'b010111101000010110110001;
#10000;
data_in <= 24'b010111101000010010101110;
#10000;
data_in <= 24'b010111011000000110101001;
#10000;
data_in <= 24'b010110010111101110011111;
#10000;
data_in <= 24'b010101100111001010010100;
#10000;
data_in <= 24'b010100100110110010001010;
#10000;
data_in <= 24'b011000111000101010110110;
#10000;
data_in <= 24'b010111111000100110110011;
#10000;
data_in <= 24'b010111111000011110110001;
#10000;
data_in <= 24'b010111111000011010101101;
#10000;
data_in <= 24'b010111011000001010101000;
#10000;
data_in <= 24'b010110010111101110011111;
#10000;
data_in <= 24'b010101010111000110010011;
#10000;
data_in <= 24'b010100010110101110001001;
#10000;
data_in <= 24'b011000001000101010110100;
#10000;
data_in <= 24'b010111101000100110110000;
#10000;
data_in <= 24'b010111101000011110101110;
#10000;
data_in <= 24'b010111101000010110101011;
#10000;
data_in <= 24'b010111001000000110100111;
#10000;
data_in <= 24'b010101110111101010011100;
#10000;
data_in <= 24'b010100010111000010001111;
#10000;
data_in <= 24'b010011100110100110000100;
#10000;
data_in <= 24'b010111111000100010101111;
#10000;
data_in <= 24'b010111011000011010101101;
#10000;
data_in <= 24'b010111101000010110101011;
#10000;
data_in <= 24'b010111001000001110101001;
#10000;
data_in <= 24'b010110100111111010100010;
#10000;
data_in <= 24'b010101000111011110011001;
#10000;
data_in <= 24'b010011100110110110001100;
#10000;
data_in <= 24'b010010110110011010000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010100010110011010000001;
#10000;
data_in <= 24'b010001010101100101101011;
#10000;
data_in <= 24'b001000010010111000111100;
#10000;
data_in <= 24'b000000000000101000010010;
#10000;
data_in <= 24'b000000000000010100001000;
#10000;
data_in <= 24'b000001110000110000001011;
#10000;
data_in <= 24'b000001100000101000000101;
#10000;
data_in <= 24'b000000110000010100000000;
#10000;
data_in <= 24'b010011110110010001111111;
#10000;
data_in <= 24'b010001100101011101101010;
#10000;
data_in <= 24'b001000100010111100111101;
#10000;
data_in <= 24'b000000000000101000010010;
#10000;
data_in <= 24'b000000000000010100001000;
#10000;
data_in <= 24'b000001100000101100001010;
#10000;
data_in <= 24'b000010010000101000000110;
#10000;
data_in <= 24'b000001100000100000000010;
#10000;
data_in <= 24'b010011100110001101111110;
#10000;
data_in <= 24'b010001010101011001101001;
#10000;
data_in <= 24'b001000100010111100111101;
#10000;
data_in <= 24'b000000010000101000010011;
#10000;
data_in <= 24'b000000000000001100000110;
#10000;
data_in <= 24'b000001000000100100001000;
#10000;
data_in <= 24'b000010010000101000001000;
#10000;
data_in <= 24'b000011000000101100000111;
#10000;
data_in <= 24'b010011010110001101111100;
#10000;
data_in <= 24'b010001010101011001101001;
#10000;
data_in <= 24'b001000100010111100111111;
#10000;
data_in <= 24'b000000010000101000010100;
#10000;
data_in <= 24'b000000000000000100000110;
#10000;
data_in <= 24'b000000110000010100000110;
#10000;
data_in <= 24'b000010010000011100000110;
#10000;
data_in <= 24'b000011010000110000001000;
#10000;
data_in <= 24'b010011000110001001111011;
#10000;
data_in <= 24'b010000100101001101100110;
#10000;
data_in <= 24'b001000000010110100111101;
#10000;
data_in <= 24'b000000010000101000010100;
#10000;
data_in <= 24'b000000000000000000001000;
#10000;
data_in <= 24'b000000010000001000000110;
#10000;
data_in <= 24'b000001110000010100000101;
#10000;
data_in <= 24'b000011010000100100001000;
#10000;
data_in <= 24'b010010000101111001110111;
#10000;
data_in <= 24'b001111010100111001100011;
#10000;
data_in <= 24'b000111000010100100111001;
#10000;
data_in <= 24'b000000000000100100010011;
#10000;
data_in <= 24'b000000000000000100001001;
#10000;
data_in <= 24'b000001000000001100000111;
#10000;
data_in <= 24'b000001100000001100000101;
#10000;
data_in <= 24'b000011000000011100001000;
#10000;
data_in <= 24'b010000110101100101110010;
#10000;
data_in <= 24'b001101100100011101011100;
#10000;
data_in <= 24'b000101100010001100110011;
#10000;
data_in <= 24'b000000000000011000010011;
#10000;
data_in <= 24'b000000010000001000001100;
#10000;
data_in <= 24'b000001110000010100001011;
#10000;
data_in <= 24'b000010000000010000001001;
#10000;
data_in <= 24'b000011000000011100001001;
#10000;
data_in <= 24'b001111100101010001101101;
#10000;
data_in <= 24'b001100010100001001010101;
#10000;
data_in <= 24'b000100010001111000101110;
#10000;
data_in <= 24'b000000000000011000010000;
#10000;
data_in <= 24'b000000100000010100001101;
#10000;
data_in <= 24'b000001110000100000001100;
#10000;
data_in <= 24'b000010010000011000001000;
#10000;
data_in <= 24'b000011010000100000001001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000111110010011000110111;
#10000;
data_in <= 24'b000110010010000000101111;
#10000;
data_in <= 24'b000010100001000100100000;
#10000;
data_in <= 24'b000010100001001000011111;
#10000;
data_in <= 24'b000101010001111000101000;
#10000;
data_in <= 24'b000011000001010100011110;
#10000;
data_in <= 24'b000000010000101000010011;
#10000;
data_in <= 24'b000010010001010100011011;
#10000;
data_in <= 24'b000110010001111000101101;
#10000;
data_in <= 24'b000110000001111100101110;
#10000;
data_in <= 24'b000011110001011000100101;
#10000;
data_in <= 24'b000010100001001000011111;
#10000;
data_in <= 24'b000011010001011000100000;
#10000;
data_in <= 24'b000011010001100000100000;
#10000;
data_in <= 24'b000010010001011000011110;
#10000;
data_in <= 24'b000010100001100000011110;
#10000;
data_in <= 24'b000101000001101100101100;
#10000;
data_in <= 24'b000101010001111000101100;
#10000;
data_in <= 24'b000101000001110100101011;
#10000;
data_in <= 24'b000010010001001000011111;
#10000;
data_in <= 24'b000000010000101100010101;
#10000;
data_in <= 24'b000010100001010100011101;
#10000;
data_in <= 24'b000011100001101100100011;
#10000;
data_in <= 24'b000001110001010000011100;
#10000;
data_in <= 24'b000111000010010000110101;
#10000;
data_in <= 24'b000100110001110100101110;
#10000;
data_in <= 24'b000101100001111000101111;
#10000;
data_in <= 24'b000010110001011000100100;
#10000;
data_in <= 24'b000000000000011100010100;
#10000;
data_in <= 24'b000000100000111000011000;
#10000;
data_in <= 24'b000010110001011100100001;
#10000;
data_in <= 24'b000000100000111100010111;
#10000;
data_in <= 24'b001010010011001101000101;
#10000;
data_in <= 24'b000101100010001100110011;
#10000;
data_in <= 24'b000101110010000100110010;
#10000;
data_in <= 24'b000101010010001000110000;
#10000;
data_in <= 24'b000010010001010000100010;
#10000;
data_in <= 24'b000001110001001100011111;
#10000;
data_in <= 24'b000011100001101000100110;
#10000;
data_in <= 24'b000010110001011100100001;
#10000;
data_in <= 24'b001010100011100001001011;
#10000;
data_in <= 24'b000111000010101000111100;
#10000;
data_in <= 24'b000110100010100000111010;
#10000;
data_in <= 24'b000111100010110100111101;
#10000;
data_in <= 24'b000110100010011100110111;
#10000;
data_in <= 24'b000101010010001000110000;
#10000;
data_in <= 24'b000110100010011100110101;
#10000;
data_in <= 24'b001000100010110100111011;
#10000;
data_in <= 24'b000111010010101101000001;
#10000;
data_in <= 24'b001000100011000101000100;
#10000;
data_in <= 24'b001000000010111101000010;
#10000;
data_in <= 24'b000111100010111000111111;
#10000;
data_in <= 24'b001000000010111001000000;
#10000;
data_in <= 24'b000111110010110100111111;
#10000;
data_in <= 24'b001001100011001001000100;
#10000;
data_in <= 24'b001100010011111001001110;
#10000;
data_in <= 24'b000010110001111000110011;
#10000;
data_in <= 24'b001000000011001101001000;
#10000;
data_in <= 24'b001000100011001101001000;
#10000;
data_in <= 24'b000101110010100000111101;
#10000;
data_in <= 24'b000110110010110001000001;
#10000;
data_in <= 24'b001000010011000001000011;
#10000;
data_in <= 24'b001001110011010101001000;
#10000;
data_in <= 24'b001101100100000101010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000001100001010000011010;
#10000;
data_in <= 24'b000001010001001000011010;
#10000;
data_in <= 24'b000010110001101000100011;
#10000;
data_in <= 24'b000101000010010000110000;
#10000;
data_in <= 24'b000100100010001100110000;
#10000;
data_in <= 24'b000010010001110000101011;
#10000;
data_in <= 24'b000101000010011000110111;
#10000;
data_in <= 24'b001001100011100101001110;
#10000;
data_in <= 24'b000000010001000100010111;
#10000;
data_in <= 24'b000000000000111000010101;
#10000;
data_in <= 24'b000001110001011000011111;
#10000;
data_in <= 24'b000101110010011100110011;
#10000;
data_in <= 24'b000111100010111000111011;
#10000;
data_in <= 24'b000101100010011100110100;
#10000;
data_in <= 24'b000101100010010100110101;
#10000;
data_in <= 24'b000110010010101000111101;
#10000;
data_in <= 24'b000011100001101100100011;
#10000;
data_in <= 24'b000001010001010100011100;
#10000;
data_in <= 24'b000001100001010100011110;
#10000;
data_in <= 24'b000100010001111100101011;
#10000;
data_in <= 24'b000110000010010100110011;
#10000;
data_in <= 24'b000100100010001000101111;
#10000;
data_in <= 24'b000100110010000000110000;
#10000;
data_in <= 24'b000101000010001100110110;
#10000;
data_in <= 24'b000010010001010100011111;
#10000;
data_in <= 24'b000001100001001000011100;
#10000;
data_in <= 24'b000010010001010100100001;
#10000;
data_in <= 24'b000011010001101100100111;
#10000;
data_in <= 24'b000100100001110100101011;
#10000;
data_in <= 24'b000011110001110000101100;
#10000;
data_in <= 24'b000100110001110100101111;
#10000;
data_in <= 24'b000101000010001000110101;
#10000;
data_in <= 24'b000000000000011100010011;
#10000;
data_in <= 24'b000000000000100100010101;
#10000;
data_in <= 24'b000001010001000100011101;
#10000;
data_in <= 24'b000100100001110100101011;
#10000;
data_in <= 24'b000111010010010100110110;
#10000;
data_in <= 24'b000110110010010100110110;
#10000;
data_in <= 24'b000101110001111000110001;
#10000;
data_in <= 24'b000011010001100000101100;
#10000;
data_in <= 24'b000110000010001100110001;
#10000;
data_in <= 24'b000011110001101000101000;
#10000;
data_in <= 24'b000010010001001000100000;
#10000;
data_in <= 24'b000011010001010100100110;
#10000;
data_in <= 24'b000110000010000000110001;
#10000;
data_in <= 24'b000111010010010100110110;
#10000;
data_in <= 24'b000100110001101000101101;
#10000;
data_in <= 24'b000000110000110100011111;
#10000;
data_in <= 24'b010000100100110001011101;
#10000;
data_in <= 24'b001101000011111001001111;
#10000;
data_in <= 24'b001000000010100000111001;
#10000;
data_in <= 24'b000011010001010000100111;
#10000;
data_in <= 24'b000010000000111000100001;
#10000;
data_in <= 24'b000010100001000000100011;
#10000;
data_in <= 24'b000010000000111000100001;
#10000;
data_in <= 24'b000000000000011100011010;
#10000;
data_in <= 24'b010001100101000101100101;
#10000;
data_in <= 24'b010010000101001001100100;
#10000;
data_in <= 24'b001110100100001101010111;
#10000;
data_in <= 24'b000111100010010100111000;
#10000;
data_in <= 24'b000001000000101100011110;
#10000;
data_in <= 24'b000000000000001000010101;
#10000;
data_in <= 24'b000000000000010000010111;
#10000;
data_in <= 24'b000000000000011100011010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101100100101101100110;
#10000;
data_in <= 24'b010000110101100001110111;
#10000;
data_in <= 24'b010010110110000001111111;
#10000;
data_in <= 24'b010010100110000110000001;
#10000;
data_in <= 24'b010010110110001110000111;
#10000;
data_in <= 24'b010010010110001110001000;
#10000;
data_in <= 24'b010011010110011110001111;
#10000;
data_in <= 24'b010110000111010010011101;
#10000;
data_in <= 24'b001010110011111101011000;
#10000;
data_in <= 24'b001110110101000001101100;
#10000;
data_in <= 24'b010001100101101101110111;
#10000;
data_in <= 24'b010010100101111101111110;
#10000;
data_in <= 24'b010011010110001110000110;
#10000;
data_in <= 24'b010010100110001010000110;
#10000;
data_in <= 24'b010011010110011110001100;
#10000;
data_in <= 24'b010110000111001010011010;
#10000;
data_in <= 24'b000111000010111001000101;
#10000;
data_in <= 24'b001011010100001001011101;
#10000;
data_in <= 24'b001111100101001101101111;
#10000;
data_in <= 24'b010001110101110001111011;
#10000;
data_in <= 24'b010011000110001010000101;
#10000;
data_in <= 24'b010010100110001010000110;
#10000;
data_in <= 24'b010010100110010010001001;
#10000;
data_in <= 24'b010101000110111010010110;
#10000;
data_in <= 24'b000100100010001000111001;
#10000;
data_in <= 24'b001001000011100001010001;
#10000;
data_in <= 24'b001110010100110001100111;
#10000;
data_in <= 24'b010001000101100101110101;
#10000;
data_in <= 24'b010011010110001010000010;
#10000;
data_in <= 24'b010010110110000110000100;
#10000;
data_in <= 24'b010010100110000110000111;
#10000;
data_in <= 24'b010100010110101110010011;
#10000;
data_in <= 24'b000011100001110000110010;
#10000;
data_in <= 24'b000111110011000101001000;
#10000;
data_in <= 24'b001100100100001101011101;
#10000;
data_in <= 24'b010000000101001101101110;
#10000;
data_in <= 24'b010010110101111101111110;
#10000;
data_in <= 24'b010011000110000010000011;
#10000;
data_in <= 24'b010010000101111110000101;
#10000;
data_in <= 24'b010011100110011110001111;
#10000;
data_in <= 24'b000011000001101000101101;
#10000;
data_in <= 24'b000110010010101000111111;
#10000;
data_in <= 24'b001010000011100001001111;
#10000;
data_in <= 24'b001101100100011101100010;
#10000;
data_in <= 24'b010001100101100001110111;
#10000;
data_in <= 24'b010010100101111101111111;
#10000;
data_in <= 24'b010010000101111010000010;
#10000;
data_in <= 24'b010010100110001110001011;
#10000;
data_in <= 24'b000010110001011100101001;
#10000;
data_in <= 24'b000100100010000100110100;
#10000;
data_in <= 24'b000110110010100101000000;
#10000;
data_in <= 24'b001010010011100001010010;
#10000;
data_in <= 24'b001111010100111101101100;
#10000;
data_in <= 24'b010001100101101001111001;
#10000;
data_in <= 24'b010001110101101101111110;
#10000;
data_in <= 24'b010010000101111110000101;
#10000;
data_in <= 24'b000010000001010000100110;
#10000;
data_in <= 24'b000011000001101000101101;
#10000;
data_in <= 24'b000100010001111100110101;
#10000;
data_in <= 24'b000111110010111001001000;
#10000;
data_in <= 24'b001110000100100101100100;
#10000;
data_in <= 24'b010000110101011101110110;
#10000;
data_in <= 24'b010001010101100101111100;
#10000;
data_in <= 24'b010001100101110110000011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011011111000110010111000;
#10000;
data_in <= 24'b100000001001110111001001;
#10000;
data_in <= 24'b100100101011001011011101;
#10000;
data_in <= 24'b100110111011110111101000;
#10000;
data_in <= 24'b100111111100001011101101;
#10000;
data_in <= 24'b100111111100011011101101;
#10000;
data_in <= 24'b101000001100011111101110;
#10000;
data_in <= 24'b100111101100010111101100;
#10000;
data_in <= 24'b011011101000100110110101;
#10000;
data_in <= 24'b011111001001110011000111;
#10000;
data_in <= 24'b100011111010111111011010;
#10000;
data_in <= 24'b100101111011101011100101;
#10000;
data_in <= 24'b100111001011111111101010;
#10000;
data_in <= 24'b100111001100001011101100;
#10000;
data_in <= 24'b100110111100001111101101;
#10000;
data_in <= 24'b100110011100000111101011;
#10000;
data_in <= 24'b011010111000011010110010;
#10000;
data_in <= 24'b011110001001100011000011;
#10000;
data_in <= 24'b100010111010101011010111;
#10000;
data_in <= 24'b100100101011010111100001;
#10000;
data_in <= 24'b100101111011101011100110;
#10000;
data_in <= 24'b100110001011110111101001;
#10000;
data_in <= 24'b100101101011110111101001;
#10000;
data_in <= 24'b100101011011110011101000;
#10000;
data_in <= 24'b011001101000001010101011;
#10000;
data_in <= 24'b011101011001001010111110;
#10000;
data_in <= 24'b100001101010010111010010;
#10000;
data_in <= 24'b100011011011000011011100;
#10000;
data_in <= 24'b100100001011010111100001;
#10000;
data_in <= 24'b100100011011100011100100;
#10000;
data_in <= 24'b100100101011100111100101;
#10000;
data_in <= 24'b100100011011100011100100;
#10000;
data_in <= 24'b011000110111110010100110;
#10000;
data_in <= 24'b011011111000110010111000;
#10000;
data_in <= 24'b100000001001111111001100;
#10000;
data_in <= 24'b100001111010101011010110;
#10000;
data_in <= 24'b100010101010111011011100;
#10000;
data_in <= 24'b100011001011001111100000;
#10000;
data_in <= 24'b100011101011010111100010;
#10000;
data_in <= 24'b100010111011010011100001;
#10000;
data_in <= 24'b010111000111010110011111;
#10000;
data_in <= 24'b011010001000010110110001;
#10000;
data_in <= 24'b011110011001100011000101;
#10000;
data_in <= 24'b100000011010010011010000;
#10000;
data_in <= 24'b100001001010100011010110;
#10000;
data_in <= 24'b100001111010111011011011;
#10000;
data_in <= 24'b100001111011000011011101;
#10000;
data_in <= 24'b100010001011000111011110;
#10000;
data_in <= 24'b010101000110110110010111;
#10000;
data_in <= 24'b011000010111111010101010;
#10000;
data_in <= 24'b011100101001000110111110;
#10000;
data_in <= 24'b011110101001110011001010;
#10000;
data_in <= 24'b011111101010001011010010;
#10000;
data_in <= 24'b100000101010100011011000;
#10000;
data_in <= 24'b100000111010101111011011;
#10000;
data_in <= 24'b100001001010110011011100;
#10000;
data_in <= 24'b010100000110100110010011;
#10000;
data_in <= 24'b010111100111100110100101;
#10000;
data_in <= 24'b011011011000110010111001;
#10000;
data_in <= 24'b011101111001100011000110;
#10000;
data_in <= 24'b011111001001110111001110;
#10000;
data_in <= 24'b100000001010010011010100;
#10000;
data_in <= 24'b100000101010100011011000;
#10000;
data_in <= 24'b100000011010100111011001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100111111100001011101101;
#10000;
data_in <= 24'b101000011100010011101111;
#10000;
data_in <= 24'b101000111100011011101110;
#10000;
data_in <= 24'b101000111100100011101110;
#10000;
data_in <= 24'b101001001100100011101100;
#10000;
data_in <= 24'b101001011100101111101101;
#10000;
data_in <= 24'b101001111100110111101111;
#10000;
data_in <= 24'b101010011100111111110001;
#10000;
data_in <= 24'b100110101011111111101011;
#10000;
data_in <= 24'b100111101100000111101101;
#10000;
data_in <= 24'b100111111100001011101101;
#10000;
data_in <= 24'b101000001100010011101100;
#10000;
data_in <= 24'b101000001100011011101001;
#10000;
data_in <= 24'b101000101100100011101010;
#10000;
data_in <= 24'b101000101100101111101100;
#10000;
data_in <= 24'b101001011100111011101110;
#10000;
data_in <= 24'b100101101011101011101000;
#10000;
data_in <= 24'b100110001011110111101001;
#10000;
data_in <= 24'b100110011011111111101001;
#10000;
data_in <= 24'b100110101100000111101000;
#10000;
data_in <= 24'b100110101100000111100111;
#10000;
data_in <= 24'b100111001100010011100111;
#10000;
data_in <= 24'b100111101100011111101000;
#10000;
data_in <= 24'b101000001100100111101010;
#10000;
data_in <= 24'b100100101011011011100100;
#10000;
data_in <= 24'b100101001011100011100110;
#10000;
data_in <= 24'b100101011011101011100110;
#10000;
data_in <= 24'b100101101011110011100110;
#10000;
data_in <= 24'b100101101011110111100100;
#10000;
data_in <= 24'b100110001011111111100101;
#10000;
data_in <= 24'b100110101100001011100101;
#10000;
data_in <= 24'b100111001100010011100111;
#10000;
data_in <= 24'b100011011011001111100011;
#10000;
data_in <= 24'b100011101011010111100010;
#10000;
data_in <= 24'b100011111011011011100010;
#10000;
data_in <= 24'b100100001011100011100010;
#10000;
data_in <= 24'b100100111011100111100011;
#10000;
data_in <= 24'b100101001011101111100010;
#10000;
data_in <= 24'b100101111011111011100101;
#10000;
data_in <= 24'b100110011100000011100110;
#10000;
data_in <= 24'b100010011010111111011111;
#10000;
data_in <= 24'b100010101011000011100000;
#10000;
data_in <= 24'b100010111011001011011111;
#10000;
data_in <= 24'b100011001011001111011111;
#10000;
data_in <= 24'b100011101011001111011111;
#10000;
data_in <= 24'b100100001011011011100000;
#10000;
data_in <= 24'b100100101011100011100010;
#10000;
data_in <= 24'b100101011011101111100101;
#10000;
data_in <= 24'b100000101010101011011010;
#10000;
data_in <= 24'b100001001010110011011100;
#10000;
data_in <= 24'b100001011010111011011011;
#10000;
data_in <= 24'b100001101011000011011011;
#10000;
data_in <= 24'b100010001010111111011011;
#10000;
data_in <= 24'b100011001011000111011101;
#10000;
data_in <= 24'b100011101011001111011111;
#10000;
data_in <= 24'b100100101011010111100001;
#10000;
data_in <= 24'b011111111010011111010111;
#10000;
data_in <= 24'b100000011010100111011001;
#10000;
data_in <= 24'b100000101010101111011000;
#10000;
data_in <= 24'b100000111010110011011001;
#10000;
data_in <= 24'b100001011010110011011001;
#10000;
data_in <= 24'b100010011010111011011010;
#10000;
data_in <= 24'b100011011011000011011100;
#10000;
data_in <= 24'b100011111011001011011110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101001111100110111110000;
#10000;
data_in <= 24'b101001101100110011101111;
#10000;
data_in <= 24'b101001001100100011110000;
#10000;
data_in <= 24'b101000001100011011110000;
#10000;
data_in <= 24'b100111101100001011110000;
#10000;
data_in <= 24'b100101111011110111101101;
#10000;
data_in <= 24'b100100001011001111100101;
#10000;
data_in <= 24'b100010001010100111100001;
#10000;
data_in <= 24'b101001011100111011101111;
#10000;
data_in <= 24'b101000101100101011101101;
#10000;
data_in <= 24'b101000001100011111101110;
#10000;
data_in <= 24'b100111101100010011101110;
#10000;
data_in <= 24'b100111001100000011101110;
#10000;
data_in <= 24'b100100111011100011101010;
#10000;
data_in <= 24'b100010001010101011100000;
#10000;
data_in <= 24'b011111101001110111011010;
#10000;
data_in <= 24'b101001101100110011101111;
#10000;
data_in <= 24'b101000101100100011101011;
#10000;
data_in <= 24'b100111101100001011101010;
#10000;
data_in <= 24'b100111011100000011101100;
#10000;
data_in <= 24'b100110101011101111101100;
#10000;
data_in <= 24'b100011011011000011100010;
#10000;
data_in <= 24'b011111101001110111010100;
#10000;
data_in <= 24'b011100101000111111001100;
#10000;
data_in <= 24'b101001001100100111101111;
#10000;
data_in <= 24'b100111101100001111101001;
#10000;
data_in <= 24'b100110101011110111101000;
#10000;
data_in <= 24'b100110101011110111101001;
#10000;
data_in <= 24'b100101101011011111101001;
#10000;
data_in <= 24'b100001111010011111011100;
#10000;
data_in <= 24'b011100111001000011001001;
#10000;
data_in <= 24'b011001011000000110111110;
#10000;
data_in <= 24'b100111111100001111101011;
#10000;
data_in <= 24'b100110011011110011100111;
#10000;
data_in <= 24'b100101111011100011100101;
#10000;
data_in <= 24'b100110001011100111100111;
#10000;
data_in <= 24'b100100011011000011100101;
#10000;
data_in <= 24'b011111101001110011010011;
#10000;
data_in <= 24'b011010011000010010111101;
#10000;
data_in <= 24'b010110110111010010110010;
#10000;
data_in <= 24'b100110111011111011101001;
#10000;
data_in <= 24'b100101011011100011100100;
#10000;
data_in <= 24'b100101001011010111100011;
#10000;
data_in <= 24'b100101001011010011100101;
#10000;
data_in <= 24'b100010111010011111011101;
#10000;
data_in <= 24'b011100111000111011000111;
#10000;
data_in <= 24'b010111000111011010110010;
#10000;
data_in <= 24'b010101000110100110100111;
#10000;
data_in <= 24'b100110001011100111100110;
#10000;
data_in <= 24'b100100111011010011100010;
#10000;
data_in <= 24'b100100111011000111100010;
#10000;
data_in <= 24'b100100011010111011100001;
#10000;
data_in <= 24'b100000111001110011010100;
#10000;
data_in <= 24'b011001110111111110111001;
#10000;
data_in <= 24'b010100000110100010100100;
#10000;
data_in <= 24'b010010110101110110011100;
#10000;
data_in <= 24'b100101101011011111100101;
#10000;
data_in <= 24'b100100101011001011100011;
#10000;
data_in <= 24'b100100101010111111100010;
#10000;
data_in <= 24'b100011101010101011100000;
#10000;
data_in <= 24'b011111011001011011001110;
#10000;
data_in <= 24'b010111100111011010110000;
#10000;
data_in <= 24'b010010010101111010011011;
#10000;
data_in <= 24'b010001000101011010010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100000001001101011100000;
#10000;
data_in <= 24'b011110011001000011011011;
#10000;
data_in <= 24'b011100011000011011010001;
#10000;
data_in <= 24'b011011011000000011001011;
#10000;
data_in <= 24'b011010000111100011000100;
#10000;
data_in <= 24'b011000100111000110111010;
#10000;
data_in <= 24'b010111010110101010110100;
#10000;
data_in <= 24'b010111000110101010110010;
#10000;
data_in <= 24'b011111001001010111011111;
#10000;
data_in <= 24'b011101101000101111011100;
#10000;
data_in <= 24'b011100001000010011010010;
#10000;
data_in <= 24'b011010110111110111001010;
#10000;
data_in <= 24'b011001000111000110111111;
#10000;
data_in <= 24'b010101010110001010101110;
#10000;
data_in <= 24'b010010110101011010100000;
#10000;
data_in <= 24'b010010000101000110011010;
#10000;
data_in <= 24'b011101001000101011010010;
#10000;
data_in <= 24'b011100001000001011001111;
#10000;
data_in <= 24'b011010000111101111000110;
#10000;
data_in <= 24'b011000000111000110111010;
#10000;
data_in <= 24'b010101000110001110101011;
#10000;
data_in <= 24'b010001010101010010011001;
#10000;
data_in <= 24'b001111010100101110001101;
#10000;
data_in <= 24'b001111010100100110001001;
#10000;
data_in <= 24'b011001010111101010111110;
#10000;
data_in <= 24'b010111110111000110111000;
#10000;
data_in <= 24'b010101100110011010101011;
#10000;
data_in <= 24'b010010010101101010011101;
#10000;
data_in <= 24'b001111110100111110010001;
#10000;
data_in <= 24'b010000000100111110001101;
#10000;
data_in <= 24'b010011100101110010010111;
#10000;
data_in <= 24'b010111100110101010100100;
#10000;
data_in <= 24'b010101000110011110101010;
#10000;
data_in <= 24'b010010110101110010011111;
#10000;
data_in <= 24'b001111010100110110001111;
#10000;
data_in <= 24'b001101000100001110000001;
#10000;
data_in <= 24'b001110000100011010000001;
#10000;
data_in <= 24'b010100000101110110010101;
#10000;
data_in <= 24'b011101101000010010111001;
#10000;
data_in <= 24'b100101111010010011011000;
#10000;
data_in <= 24'b010010010101100110011011;
#10000;
data_in <= 24'b001111100100110010001110;
#10000;
data_in <= 24'b001100010100000001111111;
#10000;
data_in <= 24'b001100110100000101111100;
#10000;
data_in <= 24'b010001100101001110001011;
#10000;
data_in <= 24'b011010110111100110101101;
#10000;
data_in <= 24'b100110101010100011011001;
#10000;
data_in <= 24'b101111001100101011111010;
#10000;
data_in <= 24'b010001000101001010010100;
#10000;
data_in <= 24'b001110100100011010001000;
#10000;
data_in <= 24'b001101010100000110000001;
#10000;
data_in <= 24'b010001110101001010001110;
#10000;
data_in <= 24'b011001110111010110101010;
#10000;
data_in <= 24'b100010101001100011001001;
#10000;
data_in <= 24'b101010011011010111100101;
#10000;
data_in <= 24'b101110101100011111110101;
#10000;
data_in <= 24'b010001000100111110010011;
#10000;
data_in <= 24'b001111000100010110001001;
#10000;
data_in <= 24'b001111100100011110001010;
#10000;
data_in <= 24'b010110110110011010100010;
#10000;
data_in <= 24'b100000111000111011000111;
#10000;
data_in <= 24'b100111101010101111011111;
#10000;
data_in <= 24'b101010001011001111100101;
#10000;
data_in <= 24'b101001011011001111100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010111010110100110101111;
#10000;
data_in <= 24'b010110010110010010101000;
#10000;
data_in <= 24'b010011100101100110011101;
#10000;
data_in <= 24'b010000010100110110001101;
#10000;
data_in <= 24'b001110100100011110000101;
#10000;
data_in <= 24'b001110110100100010000110;
#10000;
data_in <= 24'b010000010100111110001010;
#10000;
data_in <= 24'b010000110101001010010001;
#10000;
data_in <= 24'b010011010101011010011010;
#10000;
data_in <= 24'b010010110101010010010111;
#10000;
data_in <= 24'b010010000101001010010010;
#10000;
data_in <= 24'b010001110101001010010000;
#10000;
data_in <= 24'b010011000101011110010011;
#10000;
data_in <= 24'b010101100110001010011100;
#10000;
data_in <= 24'b011000000110110110100101;
#10000;
data_in <= 24'b011001010111001010110000;
#10000;
data_in <= 24'b010001110101001010010000;
#10000;
data_in <= 24'b010101100110000110011101;
#10000;
data_in <= 24'b011010110111011010110010;
#10000;
data_in <= 24'b011110011000010011000000;
#10000;
data_in <= 24'b011110111000100111000011;
#10000;
data_in <= 24'b011110101000100011000010;
#10000;
data_in <= 24'b011110111000100111000011;
#10000;
data_in <= 24'b011111101000101111001001;
#10000;
data_in <= 24'b011100000111110110110101;
#10000;
data_in <= 24'b100001011001001011001010;
#10000;
data_in <= 24'b100111111010110011100100;
#10000;
data_in <= 24'b101010111011100011110000;
#10000;
data_in <= 24'b101000001010111011101000;
#10000;
data_in <= 24'b100100011001111111011001;
#10000;
data_in <= 24'b100010011001011111010010;
#10000;
data_in <= 24'b100001111001011011010101;
#10000;
data_in <= 24'b101010111011100111101010;
#10000;
data_in <= 24'b101010001011010111101001;
#10000;
data_in <= 24'b101001101011010011101000;
#10000;
data_in <= 24'b101001101011010011101001;
#10000;
data_in <= 24'b100111101010110011100110;
#10000;
data_in <= 24'b100100101010001011011101;
#10000;
data_in <= 24'b100011011001110011011010;
#10000;
data_in <= 24'b100011001001110011011110;
#10000;
data_in <= 24'b101111111100110111111101;
#10000;
data_in <= 24'b101010001011011011100110;
#10000;
data_in <= 24'b100101011010001111010111;
#10000;
data_in <= 24'b100101011010010011011100;
#10000;
data_in <= 24'b100111001010110011100111;
#10000;
data_in <= 24'b100110001010100111101000;
#10000;
data_in <= 24'b100011011001110111100000;
#10000;
data_in <= 24'b100001001001010011011001;
#10000;
data_in <= 24'b101100011100000011101110;
#10000;
data_in <= 24'b101000011010111111011111;
#10000;
data_in <= 24'b100110001010011011011010;
#10000;
data_in <= 24'b101000001010111011101000;
#10000;
data_in <= 24'b101001011011010011110011;
#10000;
data_in <= 24'b100110101010101011101101;
#10000;
data_in <= 24'b100001101001010011011100;
#10000;
data_in <= 24'b011110001000011111010000;
#10000;
data_in <= 24'b101010001011011011100110;
#10000;
data_in <= 24'b101001011011010011100101;
#10000;
data_in <= 24'b101001111011011011101110;
#10000;
data_in <= 24'b101010111011101111110110;
#10000;
data_in <= 24'b101000011011000111110011;
#10000;
data_in <= 24'b100011001001101111100011;
#10000;
data_in <= 24'b011110111000100111010101;
#10000;
data_in <= 24'b011101001000010011010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101110100010110001101;
#10000;
data_in <= 24'b001010100011100110000010;
#10000;
data_in <= 24'b001001100011010101111101;
#10000;
data_in <= 24'b001101100100100110001100;
#10000;
data_in <= 24'b010101000110101110101001;
#10000;
data_in <= 24'b011100001000101111000100;
#10000;
data_in <= 24'b100000001001111111010100;
#10000;
data_in <= 24'b100010011010100111011010;
#10000;
data_in <= 24'b010010000101010010011100;
#10000;
data_in <= 24'b010011010101101010100110;
#10000;
data_in <= 24'b010110100110100110110010;
#10000;
data_in <= 24'b011010010111110011000000;
#10000;
data_in <= 24'b011100101000100011001001;
#10000;
data_in <= 24'b011101101001000011001100;
#10000;
data_in <= 24'b011111001001101111010000;
#10000;
data_in <= 24'b100000101010001111010100;
#10000;
data_in <= 24'b011100100111111011000110;
#10000;
data_in <= 24'b011110001000010111010001;
#10000;
data_in <= 24'b011111111000111011010111;
#10000;
data_in <= 24'b011111111001001011010110;
#10000;
data_in <= 24'b011101011000101111001100;
#10000;
data_in <= 24'b011011001000011011000010;
#10000;
data_in <= 24'b011011111000111011000011;
#10000;
data_in <= 24'b011110001001100111001010;
#10000;
data_in <= 24'b100010111001100111100001;
#10000;
data_in <= 24'b100001101001010111011110;
#10000;
data_in <= 24'b011111111000111011010110;
#10000;
data_in <= 24'b011101011000100011001100;
#10000;
data_in <= 24'b011010010111111111000000;
#10000;
data_in <= 24'b011000010111110110111001;
#10000;
data_in <= 24'b011001111000011010111011;
#10000;
data_in <= 24'b011011111001000011000001;
#10000;
data_in <= 24'b011111111000111011010011;
#10000;
data_in <= 24'b011111001000101111010011;
#10000;
data_in <= 24'b011110011000100111001110;
#10000;
data_in <= 24'b011100111000011011001001;
#10000;
data_in <= 24'b011010101000000110111111;
#10000;
data_in <= 24'b011000111000000010111001;
#10000;
data_in <= 24'b011010011000011110111110;
#10000;
data_in <= 24'b011100011001001011000100;
#10000;
data_in <= 24'b011101001000010011001001;
#10000;
data_in <= 24'b011100111000011011001010;
#10000;
data_in <= 24'b011100101000010111001000;
#10000;
data_in <= 24'b011010101000000011000001;
#10000;
data_in <= 24'b010111110111100110110101;
#10000;
data_in <= 24'b010110110111100010110001;
#10000;
data_in <= 24'b011001111000011010111101;
#10000;
data_in <= 24'b011101111001100011001010;
#10000;
data_in <= 24'b011101001000010011001001;
#10000;
data_in <= 24'b011010100111111010111111;
#10000;
data_in <= 24'b011000000111010010110101;
#10000;
data_in <= 24'b010110010111000010101110;
#10000;
data_in <= 24'b010101100111000010101100;
#10000;
data_in <= 24'b010110100111011110110000;
#10000;
data_in <= 24'b011001111000011010111101;
#10000;
data_in <= 24'b011100111001011011001000;
#10000;
data_in <= 24'b011010000111101110111110;
#10000;
data_in <= 24'b010101100110110110101011;
#10000;
data_in <= 24'b010010110110001110011111;
#10000;
data_in <= 24'b010100000110101010100110;
#10000;
data_in <= 24'b010111110111110010110101;
#10000;
data_in <= 24'b011010101000100111000000;
#10000;
data_in <= 24'b011011001000111011000011;
#10000;
data_in <= 24'b011011001000111111000001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011111101010000111001101;
#10000;
data_in <= 24'b011110001001111011001000;
#10000;
data_in <= 24'b011100101001100111000000;
#10000;
data_in <= 24'b011011011001010010111011;
#10000;
data_in <= 24'b011010111001000010110110;
#10000;
data_in <= 24'b011010001000110110110011;
#10000;
data_in <= 24'b011001101000101110110001;
#10000;
data_in <= 24'b011001001000100110101111;
#10000;
data_in <= 24'b011110111010000011001100;
#10000;
data_in <= 24'b011101111001110111000111;
#10000;
data_in <= 24'b011100011001100010111111;
#10000;
data_in <= 24'b011011001001001110111001;
#10000;
data_in <= 24'b011010101000111110110101;
#10000;
data_in <= 24'b011001111000110110110000;
#10000;
data_in <= 24'b011001001000101010101101;
#10000;
data_in <= 24'b011000101000011110101101;
#10000;
data_in <= 24'b011110001001110011001010;
#10000;
data_in <= 24'b011101001001101011000100;
#10000;
data_in <= 24'b011011111001011010111101;
#10000;
data_in <= 24'b011010101001000110110111;
#10000;
data_in <= 24'b011010001000110110110011;
#10000;
data_in <= 24'b011001011000101010110000;
#10000;
data_in <= 24'b011000101000011110101101;
#10000;
data_in <= 24'b011000001000010110101011;
#10000;
data_in <= 24'b011101011001100111000111;
#10000;
data_in <= 24'b011100101001011111000011;
#10000;
data_in <= 24'b011011011001001110111101;
#10000;
data_in <= 24'b011010001000111110110110;
#10000;
data_in <= 24'b011001111000101110110011;
#10000;
data_in <= 24'b011001001000100110101111;
#10000;
data_in <= 24'b011000001000010110101011;
#10000;
data_in <= 24'b010111101000001010101010;
#10000;
data_in <= 24'b011100101001011011000110;
#10000;
data_in <= 24'b011011111001010011000000;
#10000;
data_in <= 24'b011010111001000010111100;
#10000;
data_in <= 24'b011010001000111010111000;
#10000;
data_in <= 24'b011001111000101010110101;
#10000;
data_in <= 24'b011001001000100010110000;
#10000;
data_in <= 24'b011000101000010110101101;
#10000;
data_in <= 24'b010111111000001010101010;
#10000;
data_in <= 24'b011100001001010011000100;
#10000;
data_in <= 24'b011011101001001011000000;
#10000;
data_in <= 24'b011010111000111110111101;
#10000;
data_in <= 24'b011010011000111010111010;
#10000;
data_in <= 24'b011010011000110010111000;
#10000;
data_in <= 24'b011001101000100110110100;
#10000;
data_in <= 24'b011001001000011010110001;
#10000;
data_in <= 24'b011000011000001110101110;
#10000;
data_in <= 24'b011011111001001111000011;
#10000;
data_in <= 24'b011011011001000110111111;
#10000;
data_in <= 24'b011010111000111110111101;
#10000;
data_in <= 24'b011010101000111110111011;
#10000;
data_in <= 24'b011010101000110110111001;
#10000;
data_in <= 24'b011010001000101110110110;
#10000;
data_in <= 24'b011001101000100010110011;
#10000;
data_in <= 24'b011001001000011010110001;
#10000;
data_in <= 24'b011011111001001111000011;
#10000;
data_in <= 24'b011011011001000111000001;
#10000;
data_in <= 24'b011011001001000010111110;
#10000;
data_in <= 24'b011010111000111110111101;
#10000;
data_in <= 24'b011011001000111110111011;
#10000;
data_in <= 24'b011010101000110110111001;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011001101000100010110011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000101000011010101110;
#10000;
data_in <= 24'b011000011000010110101101;
#10000;
data_in <= 24'b010111111000010010101010;
#10000;
data_in <= 24'b010111011000000110100111;
#10000;
data_in <= 24'b010111010111111110100011;
#10000;
data_in <= 24'b010110100111101010011101;
#10000;
data_in <= 24'b010100010110111010001101;
#10000;
data_in <= 24'b010001110110001001111101;
#10000;
data_in <= 24'b011000011000010010101100;
#10000;
data_in <= 24'b011000011000010010101100;
#10000;
data_in <= 24'b010111111000001010101010;
#10000;
data_in <= 24'b010111100111111110100110;
#10000;
data_in <= 24'b010111010111110110100001;
#10000;
data_in <= 24'b010110000111011010011001;
#10000;
data_in <= 24'b010011000110100010000111;
#10000;
data_in <= 24'b010000000101101101110110;
#10000;
data_in <= 24'b011000001000001110101011;
#10000;
data_in <= 24'b011000001000001110101011;
#10000;
data_in <= 24'b011000001000000010101001;
#10000;
data_in <= 24'b010111000111110110100100;
#10000;
data_in <= 24'b010110100111101010011110;
#10000;
data_in <= 24'b010100110111000110010100;
#10000;
data_in <= 24'b010001010110000110000000;
#10000;
data_in <= 24'b001110100101001001101110;
#10000;
data_in <= 24'b010111111000000110101100;
#10000;
data_in <= 24'b011000001000001010101101;
#10000;
data_in <= 24'b011000001000000010101001;
#10000;
data_in <= 24'b010111100111110110100100;
#10000;
data_in <= 24'b010110110111100010011111;
#10000;
data_in <= 24'b010100100110111010010001;
#10000;
data_in <= 24'b010000100101101101111011;
#10000;
data_in <= 24'b001101100100110101100111;
#10000;
data_in <= 24'b011000101000001010101101;
#10000;
data_in <= 24'b011000101000001010101101;
#10000;
data_in <= 24'b011000101000000010101001;
#10000;
data_in <= 24'b010111010111110010100011;
#10000;
data_in <= 24'b010110010111011010011101;
#10000;
data_in <= 24'b010100000110101010001110;
#10000;
data_in <= 24'b010000010101100101110111;
#10000;
data_in <= 24'b001100100100011101100010;
#10000;
data_in <= 24'b011000111000001010101111;
#10000;
data_in <= 24'b011000101000001010101101;
#10000;
data_in <= 24'b011000010111111010101010;
#10000;
data_in <= 24'b010111010111101010100001;
#10000;
data_in <= 24'b010101110111001010010111;
#10000;
data_in <= 24'b010010110110011010001000;
#10000;
data_in <= 24'b001110100101001001110000;
#10000;
data_in <= 24'b001011000100001001011011;
#10000;
data_in <= 24'b011001001000001110110000;
#10000;
data_in <= 24'b011000101000001010101101;
#10000;
data_in <= 24'b010111100111101110100111;
#10000;
data_in <= 24'b010110000111010110011100;
#10000;
data_in <= 24'b010100010110101110010000;
#10000;
data_in <= 24'b010001010101111010000000;
#10000;
data_in <= 24'b001100110100100001100111;
#10000;
data_in <= 24'b001001000011100001010001;
#10000;
data_in <= 24'b011001001000001110110000;
#10000;
data_in <= 24'b011000111000000010101100;
#10000;
data_in <= 24'b010111100111101010100011;
#10000;
data_in <= 24'b010101100111000010011000;
#10000;
data_in <= 24'b010011100110011010001010;
#10000;
data_in <= 24'b010000000101011101110111;
#10000;
data_in <= 24'b001011000100000101011101;
#10000;
data_in <= 24'b000111100011000001000111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101100100110101100011;
#10000;
data_in <= 24'b001001110011100001001011;
#10000;
data_in <= 24'b000011100001101100101001;
#10000;
data_in <= 24'b000000000000011100010000;
#10000;
data_in <= 24'b000000010000010100001010;
#10000;
data_in <= 24'b000010010000101100001100;
#10000;
data_in <= 24'b000011100000110000001100;
#10000;
data_in <= 24'b000010100000100000000111;
#10000;
data_in <= 24'b001100110100101001100000;
#10000;
data_in <= 24'b001000010011001101000100;
#10000;
data_in <= 24'b000010000001010100100011;
#10000;
data_in <= 24'b000000000000010100001110;
#10000;
data_in <= 24'b000000000000010100001000;
#10000;
data_in <= 24'b000001110000100100001001;
#10000;
data_in <= 24'b000010100000101100001001;
#10000;
data_in <= 24'b000010100000100100000101;
#10000;
data_in <= 24'b001100000100010101011011;
#10000;
data_in <= 24'b000110000010101000111011;
#10000;
data_in <= 24'b000000010000111000011100;
#10000;
data_in <= 24'b000000000000010000001101;
#10000;
data_in <= 24'b000000010000011000001001;
#10000;
data_in <= 24'b000000110000011000000100;
#10000;
data_in <= 24'b000001100000011100000011;
#10000;
data_in <= 24'b000010100000101000000100;
#10000;
data_in <= 24'b001010100011111101010101;
#10000;
data_in <= 24'b000101000010010000110101;
#10000;
data_in <= 24'b000000000000101100010111;
#10000;
data_in <= 24'b000000000000011000001101;
#10000;
data_in <= 24'b000000100000011100001000;
#10000;
data_in <= 24'b000000100000010100000011;
#10000;
data_in <= 24'b000001010000011000000010;
#10000;
data_in <= 24'b000011000000110000000110;
#10000;
data_in <= 24'b001001000011011001001101;
#10000;
data_in <= 24'b000100000010000000110001;
#10000;
data_in <= 24'b000000010000110100011001;
#10000;
data_in <= 24'b000000010000100100010000;
#10000;
data_in <= 24'b000001000000100100001010;
#10000;
data_in <= 24'b000000100000010100000011;
#10000;
data_in <= 24'b000001010000011000000010;
#10000;
data_in <= 24'b000011100000111000001000;
#10000;
data_in <= 24'b000110110010111001000011;
#10000;
data_in <= 24'b000100010010000000110000;
#10000;
data_in <= 24'b000010000001001000011100;
#10000;
data_in <= 24'b000001010000110100010100;
#10000;
data_in <= 24'b000001000000100100001010;
#10000;
data_in <= 24'b000000110000011000000100;
#10000;
data_in <= 24'b000001110000100000000100;
#10000;
data_in <= 24'b000011110000111100001001;
#10000;
data_in <= 24'b000100110010010000110111;
#10000;
data_in <= 24'b000100110010000000101110;
#10000;
data_in <= 24'b000011110001100100100011;
#10000;
data_in <= 24'b000001110001000000010100;
#10000;
data_in <= 24'b000000110000100000001001;
#10000;
data_in <= 24'b000000110000011000000100;
#10000;
data_in <= 24'b000010000000100100000101;
#10000;
data_in <= 24'b000010110000110100000111;
#10000;
data_in <= 24'b000011110001111100110000;
#10000;
data_in <= 24'b000101000010000100101111;
#10000;
data_in <= 24'b000100100001110100100101;
#10000;
data_in <= 24'b000010000001000100010101;
#10000;
data_in <= 24'b000000100000011100001000;
#10000;
data_in <= 24'b000000010000011000000101;
#10000;
data_in <= 24'b000001100000101000000101;
#10000;
data_in <= 24'b000010100000110000000110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000101100010101101000001;
#10000;
data_in <= 24'b000111000011000101000111;
#10000;
data_in <= 24'b001010100011110001010011;
#10000;
data_in <= 24'b001001100011100001001111;
#10000;
data_in <= 24'b000101100010100000111111;
#10000;
data_in <= 24'b000111000010110101000010;
#10000;
data_in <= 24'b001011000011101001010000;
#10000;
data_in <= 24'b001011010011101001010000;
#10000;
data_in <= 24'b000100100010100001000001;
#10000;
data_in <= 24'b000110000010111001000111;
#10000;
data_in <= 24'b000111100011010001001101;
#10000;
data_in <= 24'b001010110011111101011000;
#10000;
data_in <= 24'b001011110100001101011100;
#10000;
data_in <= 24'b001001000011010101001111;
#10000;
data_in <= 24'b001000110011001001001100;
#10000;
data_in <= 24'b001101010100010101011100;
#10000;
data_in <= 24'b000100010010100001000010;
#10000;
data_in <= 24'b000100110010101001000100;
#10000;
data_in <= 24'b000100110010101001000100;
#10000;
data_in <= 24'b001011000100000101011100;
#10000;
data_in <= 24'b010001000101100101110100;
#10000;
data_in <= 24'b001100000100001101011110;
#10000;
data_in <= 24'b000111100011000101001100;
#10000;
data_in <= 24'b001110000100100101100100;
#10000;
data_in <= 24'b000101110011000001001010;
#10000;
data_in <= 24'b000100000010100101000011;
#10000;
data_in <= 24'b000100000010100001000100;
#10000;
data_in <= 24'b001010000011111001011010;
#10000;
data_in <= 24'b010000000101011001110010;
#10000;
data_in <= 24'b001111010101001001101110;
#10000;
data_in <= 24'b001011010100000101100000;
#10000;
data_in <= 24'b001010100011111101011011;
#10000;
data_in <= 24'b001010100100010101100000;
#10000;
data_in <= 24'b000110110011011001010001;
#10000;
data_in <= 24'b000111110011100101010111;
#10000;
data_in <= 24'b001001100011111001011100;
#10000;
data_in <= 24'b001011100100011001100100;
#10000;
data_in <= 24'b010011000110000110000000;
#10000;
data_in <= 24'b010010110110000010000000;
#10000;
data_in <= 24'b001000100011011101010110;
#10000;
data_in <= 24'b010000010101110001110111;
#10000;
data_in <= 24'b001100110100111001101001;
#10000;
data_in <= 24'b001110010101001101110001;
#10000;
data_in <= 24'b001011110100100101100111;
#10000;
data_in <= 24'b001001110011111001011110;
#10000;
data_in <= 24'b010100000110011110000111;
#10000;
data_in <= 24'b010111100111010110010101;
#10000;
data_in <= 24'b001010100100000101100001;
#10000;
data_in <= 24'b010010110110011110000101;
#10000;
data_in <= 24'b010001100110001010000000;
#10000;
data_in <= 24'b010010100110011010000101;
#10000;
data_in <= 24'b001111000101100001110111;
#10000;
data_in <= 24'b001011010100011001101000;
#10000;
data_in <= 24'b010001000101110101111111;
#10000;
data_in <= 24'b010101100110111110010001;
#10000;
data_in <= 24'b001111100101011101110111;
#10000;
data_in <= 24'b010011000110011110000010;
#10000;
data_in <= 24'b010011100110101110000110;
#10000;
data_in <= 24'b010100010110101110001001;
#10000;
data_in <= 24'b010001100110000001111110;
#10000;
data_in <= 24'b001101100100111101101111;
#10000;
data_in <= 24'b001101100100111101101111;
#10000;
data_in <= 24'b010001000101110101111101;
#10000;
data_in <= 24'b010011110110100010001000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001100010011111001010100;
#10000;
data_in <= 24'b010001100101000101100101;
#10000;
data_in <= 24'b010100010101110001110010;
#10000;
data_in <= 24'b001111110100100001011100;
#10000;
data_in <= 24'b000101110001111000110010;
#10000;
data_in <= 24'b000000000000000000010011;
#10000;
data_in <= 24'b000000000000000000010011;
#10000;
data_in <= 24'b000001100001000000100010;
#10000;
data_in <= 24'b001101010100001101011010;
#10000;
data_in <= 24'b001110010100011101011110;
#10000;
data_in <= 24'b010010110101100001101110;
#10000;
data_in <= 24'b010110000110001101111001;
#10000;
data_in <= 24'b010001010100110101100100;
#10000;
data_in <= 24'b000110010010001000110110;
#10000;
data_in <= 24'b000000000000011100011011;
#10000;
data_in <= 24'b000000000000010100010111;
#10000;
data_in <= 24'b010000100101000001101100;
#10000;
data_in <= 24'b001110100100100101100011;
#10000;
data_in <= 24'b010000000100111001100101;
#10000;
data_in <= 24'b010100010101111101110101;
#10000;
data_in <= 24'b010101100110001101111001;
#10000;
data_in <= 24'b001111100100110001011111;
#10000;
data_in <= 24'b000111100010100100111101;
#10000;
data_in <= 24'b000001010001001100100110;
#10000;
data_in <= 24'b001111000100111001101011;
#10000;
data_in <= 24'b001111000100111101101010;
#10000;
data_in <= 24'b001110010100101001100100;
#10000;
data_in <= 24'b001110010100101101100010;
#10000;
data_in <= 24'b010011000101110101110010;
#10000;
data_in <= 24'b010110000110100101111110;
#10000;
data_in <= 24'b010001010101010001100111;
#10000;
data_in <= 24'b001001000011001101000110;
#10000;
data_in <= 24'b001000110011011101010110;
#10000;
data_in <= 24'b001100010100011001100010;
#10000;
data_in <= 24'b001111000100111101101010;
#10000;
data_in <= 24'b001111110101001101101100;
#10000;
data_in <= 24'b010011100110001101111001;
#10000;
data_in <= 24'b010111010111001010000111;
#10000;
data_in <= 24'b010101000110100001111010;
#10000;
data_in <= 24'b001110110100111101100001;
#10000;
data_in <= 24'b000110110011001001010010;
#10000;
data_in <= 24'b001001000011100101011000;
#10000;
data_in <= 24'b001100010100011101100011;
#10000;
data_in <= 24'b010000000101100001110000;
#10000;
data_in <= 24'b010010000101111101110101;
#10000;
data_in <= 24'b010010010110000101110101;
#10000;
data_in <= 24'b010010110110001101110101;
#10000;
data_in <= 24'b010100010110011101111001;
#10000;
data_in <= 24'b001000100011101101011011;
#10000;
data_in <= 24'b000111100011011001010100;
#10000;
data_in <= 24'b000111010011010101010001;
#10000;
data_in <= 24'b001000100011110001010100;
#10000;
data_in <= 24'b001001110011111101010101;
#10000;
data_in <= 24'b001011010100011001011010;
#10000;
data_in <= 24'b001111100101100001101001;
#10000;
data_in <= 24'b010100010110101101111100;
#10000;
data_in <= 24'b001000100011101101011011;
#10000;
data_in <= 24'b000111010011011101010101;
#10000;
data_in <= 24'b000100010010100101000101;
#10000;
data_in <= 24'b000001000001110100110111;
#10000;
data_in <= 24'b000010000010001000111010;
#10000;
data_in <= 24'b000111100011100101001110;
#10000;
data_in <= 24'b001100100100110101100001;
#10000;
data_in <= 24'b001111010101011001101010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000001100001001000100100;
#10000;
data_in <= 24'b000001100001010000100111;
#10000;
data_in <= 24'b000100100010000000110110;
#10000;
data_in <= 24'b000111110010111101000110;
#10000;
data_in <= 24'b001010110011110001010111;
#10000;
data_in <= 24'b001111010100111101101110;
#10000;
data_in <= 24'b010010010101110001111111;
#10000;
data_in <= 24'b010001010101101010000000;
#10000;
data_in <= 24'b000100100010000000110010;
#10000;
data_in <= 24'b000011000001101100101110;
#10000;
data_in <= 24'b000100110010000100110111;
#10000;
data_in <= 24'b000110100010101001000001;
#10000;
data_in <= 24'b000111110011000001001011;
#10000;
data_in <= 24'b001011110100000101100000;
#10000;
data_in <= 24'b010000010101010001110111;
#10000;
data_in <= 24'b010001100101101110000001;
#10000;
data_in <= 24'b000011110001110100110000;
#10000;
data_in <= 24'b000010000001011100101010;
#10000;
data_in <= 24'b000011110001110100110011;
#10000;
data_in <= 24'b000110100010100101000011;
#10000;
data_in <= 24'b000111010010111001001001;
#10000;
data_in <= 24'b001010000011101001011001;
#10000;
data_in <= 24'b001110100100110101110000;
#10000;
data_in <= 24'b010000010101011001111100;
#10000;
data_in <= 24'b000010110001101000101101;
#10000;
data_in <= 24'b000000010001001000100111;
#10000;
data_in <= 24'b000010110001101100110010;
#10000;
data_in <= 24'b000111010010111001001000;
#10000;
data_in <= 24'b001001010011011101010100;
#10000;
data_in <= 24'b001010100011111001011101;
#10000;
data_in <= 24'b001101000100011101101010;
#10000;
data_in <= 24'b001101100100100101101110;
#10000;
data_in <= 24'b000111010011000001000101;
#10000;
data_in <= 24'b000011010010000000110101;
#10000;
data_in <= 24'b000011000001111000110101;
#10000;
data_in <= 24'b000110100010101101000101;
#10000;
data_in <= 24'b001001000011011001010011;
#10000;
data_in <= 24'b001011110100001001100011;
#10000;
data_in <= 24'b001110010100110001101111;
#10000;
data_in <= 24'b001110000100101101110000;
#10000;
data_in <= 24'b001110010100111001100011;
#10000;
data_in <= 24'b001001100011100001001111;
#10000;
data_in <= 24'b000101100010011101000001;
#10000;
data_in <= 24'b000011110010001000111101;
#10000;
data_in <= 24'b000101100010100001000101;
#10000;
data_in <= 24'b001011100100000101100010;
#10000;
data_in <= 24'b010010100101111010000001;
#10000;
data_in <= 24'b010101100110100110001110;
#10000;
data_in <= 24'b010011010110001001110111;
#10000;
data_in <= 24'b010000100101011101101101;
#10000;
data_in <= 24'b001011100100001001011011;
#10000;
data_in <= 24'b000100110010011001000001;
#10000;
data_in <= 24'b000010000001101000110111;
#10000;
data_in <= 24'b001000100011010101010110;
#10000;
data_in <= 24'b010011100110001010000101;
#10000;
data_in <= 24'b011001010111100010011101;
#10000;
data_in <= 24'b010110000110111010000111;
#10000;
data_in <= 24'b010110110110111110001000;
#10000;
data_in <= 24'b010011000101111101111010;
#10000;
data_in <= 24'b001000000011010101010001;
#10000;
data_in <= 24'b000000000001001100110010;
#10000;
data_in <= 24'b000100000010010101000101;
#10000;
data_in <= 24'b001111010101000001110101;
#10000;
data_in <= 24'b010101110110101010010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010001110110000010001000;
#10000;
data_in <= 24'b010101110111000010011100;
#10000;
data_in <= 24'b011001011000001010101111;
#10000;
data_in <= 24'b011011011000110010111001;
#10000;
data_in <= 24'b011100011001001111000001;
#10000;
data_in <= 24'b011101101001101011001000;
#10000;
data_in <= 24'b011110101001111011001110;
#10000;
data_in <= 24'b011110001001111011001110;
#10000;
data_in <= 24'b010001000101101010000011;
#10000;
data_in <= 24'b010100010110100110010011;
#10000;
data_in <= 24'b011000000111101110100111;
#10000;
data_in <= 24'b011010011000011010110011;
#10000;
data_in <= 24'b011011011000111010111100;
#10000;
data_in <= 24'b011100111001010111000011;
#10000;
data_in <= 24'b011101101001100011000110;
#10000;
data_in <= 24'b011101001001100011001000;
#10000;
data_in <= 24'b001111100101010001111101;
#10000;
data_in <= 24'b010010010110000110001011;
#10000;
data_in <= 24'b010110000111000110011101;
#10000;
data_in <= 24'b011000100111110110101001;
#10000;
data_in <= 24'b011010011000011010110011;
#10000;
data_in <= 24'b011011101000110110111010;
#10000;
data_in <= 24'b011100101001000110111110;
#10000;
data_in <= 24'b011100001001000110111111;
#10000;
data_in <= 24'b001111010101000101111010;
#10000;
data_in <= 24'b010001000101101010000011;
#10000;
data_in <= 24'b010100000110100010010010;
#10000;
data_in <= 24'b010111000111010110100001;
#10000;
data_in <= 24'b011001000111111110101011;
#10000;
data_in <= 24'b011010101000011110110011;
#10000;
data_in <= 24'b011011101000101110111000;
#10000;
data_in <= 24'b011011011000110010111001;
#10000;
data_in <= 24'b001111110101001101111100;
#10000;
data_in <= 24'b010000010101011110000000;
#10000;
data_in <= 24'b010010110110000110001011;
#10000;
data_in <= 24'b010101100110111010011000;
#10000;
data_in <= 24'b011000100111101010100100;
#10000;
data_in <= 24'b011010011000001010101100;
#10000;
data_in <= 24'b011011011000011010110010;
#10000;
data_in <= 24'b011011001000100110110101;
#10000;
data_in <= 24'b010000010101011001111100;
#10000;
data_in <= 24'b010000010101010101111110;
#10000;
data_in <= 24'b010001100101100110000100;
#10000;
data_in <= 24'b010100010110011110010001;
#10000;
data_in <= 24'b010111100111010010011110;
#10000;
data_in <= 24'b011001000111110110100101;
#10000;
data_in <= 24'b011010101000001010101100;
#10000;
data_in <= 24'b011010111000011110110000;
#10000;
data_in <= 24'b010001000101011101111101;
#10000;
data_in <= 24'b001111100101001101111001;
#10000;
data_in <= 24'b010000000101010001111101;
#10000;
data_in <= 24'b010010010101111110001000;
#10000;
data_in <= 24'b010101110110110110010110;
#10000;
data_in <= 24'b011000000111011110011101;
#10000;
data_in <= 24'b011001110111110110100110;
#10000;
data_in <= 24'b011010011000001110101011;
#10000;
data_in <= 24'b010001010101100001111110;
#10000;
data_in <= 24'b001111000101000001111001;
#10000;
data_in <= 24'b001110110100111101111000;
#10000;
data_in <= 24'b010001100101101010000011;
#10000;
data_in <= 24'b010101000110100010010001;
#10000;
data_in <= 24'b010111100111001110011001;
#10000;
data_in <= 24'b011001010111101010100000;
#10000;
data_in <= 24'b011001111000000010101000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011110001010000011010000;
#10000;
data_in <= 24'b011110101010001011010010;
#10000;
data_in <= 24'b011111101010010011010100;
#10000;
data_in <= 24'b011111111010011011010011;
#10000;
data_in <= 24'b100000101010011011010100;
#10000;
data_in <= 24'b100001011010100111010111;
#10000;
data_in <= 24'b100010101010110011011010;
#10000;
data_in <= 24'b100011001010111011011100;
#10000;
data_in <= 24'b011101011001101111001011;
#10000;
data_in <= 24'b011101111001110111001101;
#10000;
data_in <= 24'b011110011001111111001111;
#10000;
data_in <= 24'b011110111010000111010001;
#10000;
data_in <= 24'b011111111010001111010001;
#10000;
data_in <= 24'b100000101010011011010100;
#10000;
data_in <= 24'b100010001010101011011000;
#10000;
data_in <= 24'b100010101010110011011010;
#10000;
data_in <= 24'b011100001001010011000010;
#10000;
data_in <= 24'b011100101001011011000100;
#10000;
data_in <= 24'b011101011001100111000111;
#10000;
data_in <= 24'b011110001001110011001010;
#10000;
data_in <= 24'b011111011001111111001101;
#10000;
data_in <= 24'b100000001010001011010000;
#10000;
data_in <= 24'b100001011010010111010110;
#10000;
data_in <= 24'b100010001010100011011001;
#10000;
data_in <= 24'b011010111000111010111010;
#10000;
data_in <= 24'b011011001001000110111101;
#10000;
data_in <= 24'b011100011001001111000001;
#10000;
data_in <= 24'b011101011001011111000101;
#10000;
data_in <= 24'b011110001001101011001000;
#10000;
data_in <= 24'b011111011001111111001101;
#10000;
data_in <= 24'b100000101010001011010011;
#10000;
data_in <= 24'b100001101010011011010111;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011010101000110110111000;
#10000;
data_in <= 24'b011011111001000010111101;
#10000;
data_in <= 24'b011100101001001111000000;
#10000;
data_in <= 24'b011101101001011111000100;
#10000;
data_in <= 24'b011110101001101111001000;
#10000;
data_in <= 24'b011111111010000011001110;
#10000;
data_in <= 24'b100000101010001111010001;
#10000;
data_in <= 24'b011010101000100010110001;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011011101000111010111001;
#10000;
data_in <= 24'b011011111001000110111100;
#10000;
data_in <= 24'b011100101001001111000000;
#10000;
data_in <= 24'b011101101001011111000100;
#10000;
data_in <= 24'b011110111001110011001010;
#10000;
data_in <= 24'b011111101001111111001101;
#10000;
data_in <= 24'b011010101000011010101111;
#10000;
data_in <= 24'b011010001000100010110001;
#10000;
data_in <= 24'b011011011000101010110110;
#10000;
data_in <= 24'b011011101000111010111001;
#10000;
data_in <= 24'b011100011001000010111101;
#10000;
data_in <= 24'b011101001001001111000000;
#10000;
data_in <= 24'b011110001001011011000101;
#10000;
data_in <= 24'b011110111001100111001000;
#10000;
data_in <= 24'b011010011000010110101110;
#10000;
data_in <= 24'b011001111000011110110000;
#10000;
data_in <= 24'b011010111000100010110100;
#10000;
data_in <= 24'b011011001000110010110111;
#10000;
data_in <= 24'b011011101000111010111001;
#10000;
data_in <= 24'b011100011001000010111101;
#10000;
data_in <= 24'b011101011001010011000001;
#10000;
data_in <= 24'b011110001001011111000100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100100111011001111100100;
#10000;
data_in <= 24'b100011011010110111011110;
#10000;
data_in <= 24'b100011111010110011011111;
#10000;
data_in <= 24'b100100001010101011100000;
#10000;
data_in <= 24'b011110111001001011001010;
#10000;
data_in <= 24'b010100110110100110100011;
#10000;
data_in <= 24'b001110000100110110001010;
#10000;
data_in <= 24'b001100110100010110000100;
#10000;
data_in <= 24'b100011111010111111100000;
#10000;
data_in <= 24'b100011001010100111011100;
#10000;
data_in <= 24'b100011011010100111011111;
#10000;
data_in <= 24'b100010111010010111011011;
#10000;
data_in <= 24'b011100111000101011000010;
#10000;
data_in <= 24'b010010110110000110011011;
#10000;
data_in <= 24'b001100000100011010000000;
#10000;
data_in <= 24'b001010110011110101111100;
#10000;
data_in <= 24'b100011001010100111011100;
#10000;
data_in <= 24'b100011001010100111011100;
#10000;
data_in <= 24'b100011111010101111100001;
#10000;
data_in <= 24'b100010001010010011011010;
#10000;
data_in <= 24'b011011001000010110111101;
#10000;
data_in <= 24'b010000010101101010010010;
#10000;
data_in <= 24'b001000010011101001110010;
#10000;
data_in <= 24'b000110010010111001101011;
#10000;
data_in <= 24'b100001011010001011010101;
#10000;
data_in <= 24'b100010101010011111011010;
#10000;
data_in <= 24'b100011101010101011100000;
#10000;
data_in <= 24'b100001011010000111010111;
#10000;
data_in <= 24'b011010011000001010111010;
#10000;
data_in <= 24'b001111100101011110001111;
#10000;
data_in <= 24'b000111010011011001101110;
#10000;
data_in <= 24'b000100100010011101100100;
#10000;
data_in <= 24'b100000011001111111010000;
#10000;
data_in <= 24'b100001011010001111010100;
#10000;
data_in <= 24'b100001111010010011010111;
#10000;
data_in <= 24'b011111101001101111001110;
#10000;
data_in <= 24'b011010001000010010111010;
#10000;
data_in <= 24'b010011000110100010011110;
#10000;
data_in <= 24'b001101110101001110001001;
#10000;
data_in <= 24'b001011110100011110000001;
#10000;
data_in <= 24'b100000111010000111010010;
#10000;
data_in <= 24'b100001011010001111010100;
#10000;
data_in <= 24'b100000111010000011010011;
#10000;
data_in <= 24'b011111001001100111001100;
#10000;
data_in <= 24'b011100111000111111000101;
#10000;
data_in <= 24'b011011011000100110111111;
#10000;
data_in <= 24'b011010011000010110111011;
#10000;
data_in <= 24'b011001101000000110111001;
#10000;
data_in <= 24'b100000001001111011001111;
#10000;
data_in <= 24'b100000101010000011010001;
#10000;
data_in <= 24'b011111111001111111010000;
#10000;
data_in <= 24'b011111001001110011001101;
#10000;
data_in <= 24'b011111011001110011001111;
#10000;
data_in <= 24'b100000011010000011010011;
#10000;
data_in <= 24'b100000101010000111010100;
#10000;
data_in <= 24'b100000011001110111010011;
#10000;
data_in <= 24'b011101011001010011000001;
#10000;
data_in <= 24'b011110101001100111000110;
#10000;
data_in <= 24'b011110101001101111001000;
#10000;
data_in <= 24'b011110111001110011001001;
#10000;
data_in <= 24'b011111101001111111001101;
#10000;
data_in <= 24'b100000101010001111010001;
#10000;
data_in <= 24'b011111101001111111001101;
#10000;
data_in <= 24'b011101011001011011000100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010000010100101110010001;
#10000;
data_in <= 24'b001011000011010001111010;
#10000;
data_in <= 24'b001110010100000010000101;
#10000;
data_in <= 24'b011100010111101010111010;
#10000;
data_in <= 24'b100111011010011111100011;
#10000;
data_in <= 24'b101000001010101111100100;
#10000;
data_in <= 24'b100110011010010111011011;
#10000;
data_in <= 24'b100111011010101011011110;
#10000;
data_in <= 24'b001011100011101010000000;
#10000;
data_in <= 24'b001100000011011110000000;
#10000;
data_in <= 24'b010001100100111010010100;
#10000;
data_in <= 24'b011100110111110010111111;
#10000;
data_in <= 24'b100101001001110111011100;
#10000;
data_in <= 24'b100110011010001111011111;
#10000;
data_in <= 24'b100111001010011111100001;
#10000;
data_in <= 24'b101001001011000111101001;
#10000;
data_in <= 24'b000100100010000101100110;
#10000;
data_in <= 24'b001101000011110110000110;
#10000;
data_in <= 24'b011000010110101110110001;
#10000;
data_in <= 24'b100001001000111111010011;
#10000;
data_in <= 24'b100101011001111011100001;
#10000;
data_in <= 24'b100101101010000011100000;
#10000;
data_in <= 24'b100101101010000111011111;
#10000;
data_in <= 24'b100110011010010011100010;
#10000;
data_in <= 24'b001000110011010001110111;
#10000;
data_in <= 24'b010011100101110010100100;
#10000;
data_in <= 24'b011111001000100011001110;
#10000;
data_in <= 24'b100100001001110111100001;
#10000;
data_in <= 24'b100100011001111011100010;
#10000;
data_in <= 24'b100100001001110011011110;
#10000;
data_in <= 24'b100010111001011111011001;
#10000;
data_in <= 24'b100001011001000111010001;
#10000;
data_in <= 24'b010110110110111110110000;
#10000;
data_in <= 24'b011101011000011011001001;
#10000;
data_in <= 24'b100001101001011011011001;
#10000;
data_in <= 24'b100000101001001011010101;
#10000;
data_in <= 24'b011111001000110011001111;
#10000;
data_in <= 24'b011111011000101011001110;
#10000;
data_in <= 24'b011110011000011011001010;
#10000;
data_in <= 24'b011011110111110110111111;
#10000;
data_in <= 24'b011101101000111011001010;
#10000;
data_in <= 24'b011111011001001011010000;
#10000;
data_in <= 24'b011110011000110111001110;
#10000;
data_in <= 24'b011011111000000111000010;
#10000;
data_in <= 24'b011001010111011010111001;
#10000;
data_in <= 24'b011000000111000010110011;
#10000;
data_in <= 24'b010101100110011010101001;
#10000;
data_in <= 24'b010010100101101010011100;
#10000;
data_in <= 24'b011010111000011010111110;
#10000;
data_in <= 24'b011010001000000010111010;
#10000;
data_in <= 24'b011000000111100010110100;
#10000;
data_in <= 24'b010110110111000010101110;
#10000;
data_in <= 24'b010100100110011010100111;
#10000;
data_in <= 24'b010010010101101010011101;
#10000;
data_in <= 24'b001111110101000010010011;
#10000;
data_in <= 24'b001110010100101110001100;
#10000;
data_in <= 24'b011001111000010010110111;
#10000;
data_in <= 24'b010110010111010110101011;
#10000;
data_in <= 24'b010011000110011110011111;
#10000;
data_in <= 24'b010010000110000010011010;
#10000;
data_in <= 24'b010000100101101010010110;
#10000;
data_in <= 24'b001111000101001110010001;
#10000;
data_in <= 24'b010000010101011010010100;
#10000;
data_in <= 24'b010010010101111010011011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101110101100011011111100;
#10000;
data_in <= 24'b101011011011101011110010;
#10000;
data_in <= 24'b100110101010100011100011;
#10000;
data_in <= 24'b100011101001110111011100;
#10000;
data_in <= 24'b100010101001100111011110;
#10000;
data_in <= 24'b100000111001001011011011;
#10000;
data_in <= 24'b011100000111110111001011;
#10000;
data_in <= 24'b010110110110101110110111;
#10000;
data_in <= 24'b101000011010110111100111;
#10000;
data_in <= 24'b100110101010100011100011;
#10000;
data_in <= 24'b100011111001111011011100;
#10000;
data_in <= 24'b100001001001010011010110;
#10000;
data_in <= 24'b011101101000011011001011;
#10000;
data_in <= 24'b011000110111010010111101;
#10000;
data_in <= 24'b010100100110001010101111;
#10000;
data_in <= 24'b010001000101100010011111;
#10000;
data_in <= 24'b100011101001100111010111;
#10000;
data_in <= 24'b100001101001001111010001;
#10000;
data_in <= 24'b011111001000101111001010;
#10000;
data_in <= 24'b011011100111111011000000;
#10000;
data_in <= 24'b010110000110100110101100;
#10000;
data_in <= 24'b010000000101001110010111;
#10000;
data_in <= 24'b001110000100100110010010;
#10000;
data_in <= 24'b001110010100111110010001;
#10000;
data_in <= 24'b011111011000100111001001;
#10000;
data_in <= 24'b011010110111101010111001;
#10000;
data_in <= 24'b010110010110101010101001;
#10000;
data_in <= 24'b010011000101111010011101;
#10000;
data_in <= 24'b001111000101000110001111;
#10000;
data_in <= 24'b001100100100011110000101;
#10000;
data_in <= 24'b001110010100111110010000;
#10000;
data_in <= 24'b010010100110001010011100;
#10000;
data_in <= 24'b010111000110101110101010;
#10000;
data_in <= 24'b010001010101011110010100;
#10000;
data_in <= 24'b001101000100011010000011;
#10000;
data_in <= 24'b001100110100011110000000;
#10000;
data_in <= 24'b001110010101000010001000;
#10000;
data_in <= 24'b010001000101110010010010;
#10000;
data_in <= 24'b010110000111001110100110;
#10000;
data_in <= 24'b011011101000101010111001;
#10000;
data_in <= 24'b001110010100101010001001;
#10000;
data_in <= 24'b001011100100000001111101;
#10000;
data_in <= 24'b001010100011111001110111;
#10000;
data_in <= 24'b001110100101000010000100;
#10000;
data_in <= 24'b010100010110101110011010;
#10000;
data_in <= 24'b011010001000010110110010;
#10000;
data_in <= 24'b011111101001110011000101;
#10000;
data_in <= 24'b100011011010111011010101;
#10000;
data_in <= 24'b001110010100101110001010;
#10000;
data_in <= 24'b001111110101001110001101;
#10000;
data_in <= 24'b010011010110001010011001;
#10000;
data_in <= 24'b011000100111100110101001;
#10000;
data_in <= 24'b011110001001010010111101;
#10000;
data_in <= 24'b100011001010110011010000;
#10000;
data_in <= 24'b100111001011110111011110;
#10000;
data_in <= 24'b101000101100011011100100;
#10000;
data_in <= 24'b010011110110010110011111;
#10000;
data_in <= 24'b011000000111100010101110;
#10000;
data_in <= 24'b011101011000111011000000;
#10000;
data_in <= 24'b100001101010000111001101;
#10000;
data_in <= 24'b100101001011000111010110;
#10000;
data_in <= 24'b101000011100001011100011;
#10000;
data_in <= 24'b101010111100110111101010;
#10000;
data_in <= 24'b101011011101001011101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010010100101111110011101;
#10000;
data_in <= 24'b010000100101101110010011;
#10000;
data_in <= 24'b010001100101111110010111;
#10000;
data_in <= 24'b010110000111001110101011;
#10000;
data_in <= 24'b011011001000101011000001;
#10000;
data_in <= 24'b011101011001010111001010;
#10000;
data_in <= 24'b011101001001011011001011;
#10000;
data_in <= 24'b011100111001011011001000;
#10000;
data_in <= 24'b010000010101100110010011;
#10000;
data_in <= 24'b010000110110000010010011;
#10000;
data_in <= 24'b010100010110111010100001;
#10000;
data_in <= 24'b011001001000001110110110;
#10000;
data_in <= 24'b011100111001010011000110;
#10000;
data_in <= 24'b011101111001101011001100;
#10000;
data_in <= 24'b011110011001110011001110;
#10000;
data_in <= 24'b011110101001111011001110;
#10000;
data_in <= 24'b010001100110000010010110;
#10000;
data_in <= 24'b010100100111000110011110;
#10000;
data_in <= 24'b011010001000011010110101;
#10000;
data_in <= 24'b011110001001100111000111;
#10000;
data_in <= 24'b011111111010000011010001;
#10000;
data_in <= 24'b011111101010001011010010;
#10000;
data_in <= 24'b011111111010001111010011;
#10000;
data_in <= 24'b100000001010011111010100;
#10000;
data_in <= 24'b010111100111110010101011;
#10000;
data_in <= 24'b011010111000111010110110;
#10000;
data_in <= 24'b011111101010000011001011;
#10000;
data_in <= 24'b100010011010110011010111;
#10000;
data_in <= 24'b100010001010110111011001;
#10000;
data_in <= 24'b100001011010101011010110;
#10000;
data_in <= 24'b100000111010101011010110;
#10000;
data_in <= 24'b100001011010110011011001;
#10000;
data_in <= 24'b011111111010000011000111;
#10000;
data_in <= 24'b100001011010100111001101;
#10000;
data_in <= 24'b100011011011000111010111;
#10000;
data_in <= 24'b100100011011011011011100;
#10000;
data_in <= 24'b100100001011011111011110;
#10000;
data_in <= 24'b100011101011010011011110;
#10000;
data_in <= 24'b100010101011001011011100;
#10000;
data_in <= 24'b100010001010111111011011;
#10000;
data_in <= 24'b100101111011110011011110;
#10000;
data_in <= 24'b100101111011111011011110;
#10000;
data_in <= 24'b100101111011110111011111;
#10000;
data_in <= 24'b100101011011110111100000;
#10000;
data_in <= 24'b100101111011111011100100;
#10000;
data_in <= 24'b100101111011111011100101;
#10000;
data_in <= 24'b100100011011101011100001;
#10000;
data_in <= 24'b100010111011001111011101;
#10000;
data_in <= 24'b101010011100111111101101;
#10000;
data_in <= 24'b101010001101000011101101;
#10000;
data_in <= 24'b101001011100110111101010;
#10000;
data_in <= 24'b101000011100101011101010;
#10000;
data_in <= 24'b101000011100100111101100;
#10000;
data_in <= 24'b100111101100100011101101;
#10000;
data_in <= 24'b100101011011111011100101;
#10000;
data_in <= 24'b100010111011010011011011;
#10000;
data_in <= 24'b101101101101101111110101;
#10000;
data_in <= 24'b101101101101111011110111;
#10000;
data_in <= 24'b101101001101101111110111;
#10000;
data_in <= 24'b101011101101011011110011;
#10000;
data_in <= 24'b101010101101001111110100;
#10000;
data_in <= 24'b101001011100110011110010;
#10000;
data_in <= 24'b100101111100000011100111;
#10000;
data_in <= 24'b100010101011001011011100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011100101001100011001000;
#10000;
data_in <= 24'b011011111001010111000101;
#10000;
data_in <= 24'b011011101001001011000000;
#10000;
data_in <= 24'b011010111000111110111101;
#10000;
data_in <= 24'b011010111000111010111010;
#10000;
data_in <= 24'b011010011000110010111000;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011001101000100010110011;
#10000;
data_in <= 24'b011101001001101011001010;
#10000;
data_in <= 24'b011100101001100111000110;
#10000;
data_in <= 24'b011100101001011011000100;
#10000;
data_in <= 24'b011011111001010011000000;
#10000;
data_in <= 24'b011011111001001010111110;
#10000;
data_in <= 24'b011010111000111010111001;
#10000;
data_in <= 24'b011001101000100010110011;
#10000;
data_in <= 24'b011000111000001110101110;
#10000;
data_in <= 24'b011110001001111111001100;
#10000;
data_in <= 24'b011101101001110111001010;
#10000;
data_in <= 24'b011101101001101011001000;
#10000;
data_in <= 24'b011101011001101011000110;
#10000;
data_in <= 24'b011100111001011011000010;
#10000;
data_in <= 24'b011011001000111110111010;
#10000;
data_in <= 24'b011001001000011010110001;
#10000;
data_in <= 24'b010111110111111110101000;
#10000;
data_in <= 24'b011111011010010011010001;
#10000;
data_in <= 24'b011110101010000111001101;
#10000;
data_in <= 24'b011110011001111011001010;
#10000;
data_in <= 24'b011101111001110111000111;
#10000;
data_in <= 24'b011101011001100011000011;
#10000;
data_in <= 24'b011011101001001010111010;
#10000;
data_in <= 24'b011001001000011110101111;
#10000;
data_in <= 24'b010111100111111110100110;
#10000;
data_in <= 24'b100000011010100011010100;
#10000;
data_in <= 24'b011111011010010011010000;
#10000;
data_in <= 24'b011110101001111111001011;
#10000;
data_in <= 24'b011101111001110111000111;
#10000;
data_in <= 24'b011101011001100011000011;
#10000;
data_in <= 24'b011011111001001010111010;
#10000;
data_in <= 24'b011001111000011110110000;
#10000;
data_in <= 24'b010111100111111110100110;
#10000;
data_in <= 24'b100001001010101111010111;
#10000;
data_in <= 24'b011111111010011111010001;
#10000;
data_in <= 24'b011110101010000011001010;
#10000;
data_in <= 24'b011101111001111011000101;
#10000;
data_in <= 24'b011101101001100111000001;
#10000;
data_in <= 24'b011011111001001110111001;
#10000;
data_in <= 24'b011001011000011010101101;
#10000;
data_in <= 24'b010111010111110110100001;
#10000;
data_in <= 24'b100001011010110111010111;
#10000;
data_in <= 24'b100000001010100011010010;
#10000;
data_in <= 24'b011111001010001011001100;
#10000;
data_in <= 24'b011110011010000011000111;
#10000;
data_in <= 24'b011101111001101011000010;
#10000;
data_in <= 24'b011011011001000110110111;
#10000;
data_in <= 24'b011000001000000110101000;
#10000;
data_in <= 24'b010101100111011010011001;
#10000;
data_in <= 24'b100001011010110011011000;
#10000;
data_in <= 24'b100000001010011111010011;
#10000;
data_in <= 24'b011111101010010011001110;
#10000;
data_in <= 24'b011111011010000011001011;
#10000;
data_in <= 24'b011110011001110011000100;
#10000;
data_in <= 24'b011011101000111110110110;
#10000;
data_in <= 24'b010110110111110110100001;
#10000;
data_in <= 24'b010011110110111110010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011000101000001010101101;
#10000;
data_in <= 24'b011000100111111110101011;
#10000;
data_in <= 24'b010111000111100010100001;
#10000;
data_in <= 24'b010100000110101110010000;
#10000;
data_in <= 24'b010001000101110101111111;
#10000;
data_in <= 24'b001101100100101101101010;
#10000;
data_in <= 24'b001000100011010101010000;
#10000;
data_in <= 24'b000100110010010000111001;
#10000;
data_in <= 24'b011000100111111110101011;
#10000;
data_in <= 24'b011000100111111010100111;
#10000;
data_in <= 24'b010110100111010010011100;
#10000;
data_in <= 24'b010011000110011010001010;
#10000;
data_in <= 24'b001111110101011001110110;
#10000;
data_in <= 24'b001011100100010001100000;
#10000;
data_in <= 24'b000111100010111101001001;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b010111110111110110100110;
#10000;
data_in <= 24'b010111100111101110100010;
#10000;
data_in <= 24'b010101100111001010010101;
#10000;
data_in <= 24'b010001110110000010000010;
#10000;
data_in <= 24'b001101110100110001101011;
#10000;
data_in <= 24'b001001000011100101010100;
#10000;
data_in <= 24'b000101110010011100111110;
#10000;
data_in <= 24'b000011010001101100101101;
#10000;
data_in <= 24'b010111000111101110100010;
#10000;
data_in <= 24'b010110110111011010011011;
#10000;
data_in <= 24'b010100000110101110001101;
#10000;
data_in <= 24'b001111110101100001111000;
#10000;
data_in <= 24'b001011010100001101011111;
#10000;
data_in <= 24'b000111000011000001001001;
#10000;
data_in <= 24'b000100010010001000110111;
#10000;
data_in <= 24'b000010110001100100101011;
#10000;
data_in <= 24'b010110000111100010011011;
#10000;
data_in <= 24'b010101000111000010010010;
#10000;
data_in <= 24'b010001110110001110000010;
#10000;
data_in <= 24'b001110010101000101101111;
#10000;
data_in <= 24'b001001100011101101010110;
#10000;
data_in <= 24'b000101110010100101000000;
#10000;
data_in <= 24'b000011110001111000110001;
#10000;
data_in <= 24'b000011010001101000101010;
#10000;
data_in <= 24'b010100110111001010010011;
#10000;
data_in <= 24'b010010010110011010000101;
#10000;
data_in <= 24'b001110100101011001110100;
#10000;
data_in <= 24'b001011010100010101100001;
#10000;
data_in <= 24'b000111100011010001001101;
#10000;
data_in <= 24'b000100100010010100111010;
#10000;
data_in <= 24'b000011010001101100101110;
#10000;
data_in <= 24'b000011100001100000101001;
#10000;
data_in <= 24'b010010100110100110001000;
#10000;
data_in <= 24'b001111010101101101111000;
#10000;
data_in <= 24'b001011000100100101100100;
#10000;
data_in <= 24'b001000010011101001010100;
#10000;
data_in <= 24'b000110000010110101000011;
#10000;
data_in <= 24'b000011110010000000110011;
#10000;
data_in <= 24'b000011000001100000101010;
#10000;
data_in <= 24'b000011000001011000100111;
#10000;
data_in <= 24'b010001100110001010000001;
#10000;
data_in <= 24'b001101110101001001101101;
#10000;
data_in <= 24'b001001100011111101011001;
#10000;
data_in <= 24'b000111000011001001001011;
#10000;
data_in <= 24'b000101010010011100111110;
#10000;
data_in <= 24'b000011010001110000101111;
#10000;
data_in <= 24'b000010010001010100100111;
#10000;
data_in <= 24'b000011000001010000100101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000010110001100100101011;
#10000;
data_in <= 24'b000101000010000000101100;
#10000;
data_in <= 24'b000101100001111100101000;
#10000;
data_in <= 24'b000011110001010100011010;
#10000;
data_in <= 24'b000001010000101000001101;
#10000;
data_in <= 24'b000000010000011000000101;
#10000;
data_in <= 24'b000001100000100100000111;
#10000;
data_in <= 24'b000010010000110100001000;
#10000;
data_in <= 24'b000011100001101100101011;
#10000;
data_in <= 24'b000101000001110100101010;
#10000;
data_in <= 24'b000101110001111000100111;
#10000;
data_in <= 24'b000100100001100000011111;
#10000;
data_in <= 24'b000010010000111000010001;
#10000;
data_in <= 24'b000000010000010100000110;
#10000;
data_in <= 24'b000000110000010100000101;
#10000;
data_in <= 24'b000001110000100100001001;
#10000;
data_in <= 24'b000100000001101100101001;
#10000;
data_in <= 24'b000100010001101000100111;
#10000;
data_in <= 24'b000101010001110000100101;
#10000;
data_in <= 24'b000101110001110100100100;
#10000;
data_in <= 24'b000011110001001100011000;
#10000;
data_in <= 24'b000000110000011000001010;
#10000;
data_in <= 24'b000000010000001000000110;
#10000;
data_in <= 24'b000001000000011000000111;
#10000;
data_in <= 24'b000100000001101100101001;
#10000;
data_in <= 24'b000100000001100000100101;
#10000;
data_in <= 24'b000101100001101000100101;
#10000;
data_in <= 24'b000111000001111000101000;
#10000;
data_in <= 24'b000101100001100000100000;
#10000;
data_in <= 24'b000001110000101000001111;
#10000;
data_in <= 24'b000000010000000100000111;
#10000;
data_in <= 24'b000000100000001000001000;
#10000;
data_in <= 24'b000100010001101000101000;
#10000;
data_in <= 24'b000011110001011100100100;
#10000;
data_in <= 24'b000101100001101000100101;
#10000;
data_in <= 24'b000111010001111100101001;
#10000;
data_in <= 24'b000110110001110000100110;
#10000;
data_in <= 24'b000011100000111100011001;
#10000;
data_in <= 24'b000000110000010000001110;
#10000;
data_in <= 24'b000000000000000100001011;
#10000;
data_in <= 24'b000100000001011100100110;
#10000;
data_in <= 24'b000100100001100000100101;
#10000;
data_in <= 24'b000101100001101000100101;
#10000;
data_in <= 24'b000110110001110100101000;
#10000;
data_in <= 24'b000111010001110100101001;
#10000;
data_in <= 24'b000101100001011000100010;
#10000;
data_in <= 24'b000010110000101100010111;
#10000;
data_in <= 24'b000000100000001000001110;
#10000;
data_in <= 24'b000011100001010100100100;
#10000;
data_in <= 24'b000101000001101000100111;
#10000;
data_in <= 24'b000101100001100100100111;
#10000;
data_in <= 24'b000110000001100100100111;
#10000;
data_in <= 24'b000111010001110100101011;
#10000;
data_in <= 24'b000111100001111000101100;
#10000;
data_in <= 24'b000100110001001100100001;
#10000;
data_in <= 24'b000001000000010000010010;
#10000;
data_in <= 24'b000011010001010000100011;
#10000;
data_in <= 24'b000101010001101100101000;
#10000;
data_in <= 24'b000101110001101000101000;
#10000;
data_in <= 24'b000100110001011000100100;
#10000;
data_in <= 24'b000110110001110000101010;
#10000;
data_in <= 24'b001000100010001100110001;
#10000;
data_in <= 24'b000110000001100000101000;
#10000;
data_in <= 24'b000001010000010100010101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001110010101001101101011;
#10000;
data_in <= 24'b001110100101011001101110;
#10000;
data_in <= 24'b010000100101101101110101;
#10000;
data_in <= 24'b010011000110010101111111;
#10000;
data_in <= 24'b010101100110111010001010;
#10000;
data_in <= 24'b010101110110111110001101;
#10000;
data_in <= 24'b010011100110011010000100;
#10000;
data_in <= 24'b010000110101101001111010;
#10000;
data_in <= 24'b000111110011011101001101;
#10000;
data_in <= 24'b001001100011111001010100;
#10000;
data_in <= 24'b001100110100101101100001;
#10000;
data_in <= 24'b010001100101111001110110;
#10000;
data_in <= 24'b010101110110111010001000;
#10000;
data_in <= 24'b010111010111001110001111;
#10000;
data_in <= 24'b010100110110100110000101;
#10000;
data_in <= 24'b010001100101101101111010;
#10000;
data_in <= 24'b000011000010010000111000;
#10000;
data_in <= 24'b000101110010111101000011;
#10000;
data_in <= 24'b001010000100000001010100;
#10000;
data_in <= 24'b001110110101001001101000;
#10000;
data_in <= 24'b010011000110001001111011;
#10000;
data_in <= 24'b010011110110010001111111;
#10000;
data_in <= 24'b010000010101011001110001;
#10000;
data_in <= 24'b001100000100010101100001;
#10000;
data_in <= 24'b000001100001101000101011;
#10000;
data_in <= 24'b000101100010101000111011;
#10000;
data_in <= 24'b001010000011110001001110;
#10000;
data_in <= 24'b001100110100011001011011;
#10000;
data_in <= 24'b001110000100101001100001;
#10000;
data_in <= 24'b001101010100011101011110;
#10000;
data_in <= 24'b001001100011011101010001;
#10000;
data_in <= 24'b000101100010011101000001;
#10000;
data_in <= 24'b000000000000111100011111;
#10000;
data_in <= 24'b000101010010010100110101;
#10000;
data_in <= 24'b001010000011100001001001;
#10000;
data_in <= 24'b001010100011101001001011;
#10000;
data_in <= 24'b001001100011010101001000;
#10000;
data_in <= 24'b001000100011000001000110;
#10000;
data_in <= 24'b000110110010100101000000;
#10000;
data_in <= 24'b000100110010000100111000;
#10000;
data_in <= 24'b000000000000110100011001;
#10000;
data_in <= 24'b000101110010010000110010;
#10000;
data_in <= 24'b001010010011011001000100;
#10000;
data_in <= 24'b001001000011000101000001;
#10000;
data_in <= 24'b000110010010010100110111;
#10000;
data_in <= 24'b000101100010000100110101;
#10000;
data_in <= 24'b000101110010001000110110;
#10000;
data_in <= 24'b000101010010000000110110;
#10000;
data_in <= 24'b000000110000111100011001;
#10000;
data_in <= 24'b000110100010011000110000;
#10000;
data_in <= 24'b001010000011010001000000;
#10000;
data_in <= 24'b000111100010100100110111;
#10000;
data_in <= 24'b000100010001110000101010;
#10000;
data_in <= 24'b000100000001101000101011;
#10000;
data_in <= 24'b000100110001110100101111;
#10000;
data_in <= 24'b000100100001101100101111;
#10000;
data_in <= 24'b000000100000110100010101;
#10000;
data_in <= 24'b000101110010001000101010;
#10000;
data_in <= 24'b001000100010110000110110;
#10000;
data_in <= 24'b000110010010001000101111;
#10000;
data_in <= 24'b000011100001011100100101;
#10000;
data_in <= 24'b000100000001100100100111;
#10000;
data_in <= 24'b000100110001101100101100;
#10000;
data_in <= 24'b000100100001100100101100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010000000101011101110111;
#10000;
data_in <= 24'b001001110011111001011110;
#10000;
data_in <= 24'b000011100010011001000100;
#10000;
data_in <= 24'b000001010001110100111001;
#10000;
data_in <= 24'b000000100001101000110110;
#10000;
data_in <= 24'b000001010001111000111000;
#10000;
data_in <= 24'b000101100011000001001000;
#10000;
data_in <= 24'b001011010100010101011101;
#10000;
data_in <= 24'b001111010101001001110001;
#10000;
data_in <= 24'b001010000011110101011100;
#10000;
data_in <= 24'b000101010010101001001001;
#10000;
data_in <= 24'b000100000010011001000010;
#10000;
data_in <= 24'b000011010010001100111111;
#10000;
data_in <= 24'b000010110010001000111100;
#10000;
data_in <= 24'b000100110010101001000100;
#10000;
data_in <= 24'b001000000011011101010001;
#10000;
data_in <= 24'b001100100100011101100011;
#10000;
data_in <= 24'b001000110011100001010100;
#10000;
data_in <= 24'b000110110011000001001100;
#10000;
data_in <= 24'b000111100011001101001110;
#10000;
data_in <= 24'b000111100011001101001110;
#10000;
data_in <= 24'b000101100010110001000101;
#10000;
data_in <= 24'b000100010010011101000000;
#10000;
data_in <= 24'b000101100010101001000011;
#10000;
data_in <= 24'b001000110011010001001111;
#10000;
data_in <= 24'b000111010010111001001001;
#10000;
data_in <= 24'b001000000011000101001100;
#10000;
data_in <= 24'b001011010011111001011000;
#10000;
data_in <= 24'b001100100100001101011101;
#10000;
data_in <= 24'b001010000011101001010001;
#10000;
data_in <= 24'b000110110010110101000100;
#10000;
data_in <= 24'b000101000010011000111101;
#10000;
data_in <= 24'b000101000010000100111011;
#10000;
data_in <= 24'b000101010010001100111010;
#10000;
data_in <= 24'b001000000010111001000101;
#10000;
data_in <= 24'b001100110100000101010111;
#10000;
data_in <= 24'b001111010100101101100001;
#10000;
data_in <= 24'b001101010100010001010111;
#10000;
data_in <= 24'b001001100011010101001000;
#10000;
data_in <= 24'b000110110010110000111111;
#10000;
data_in <= 24'b000011100001100100101111;
#10000;
data_in <= 24'b000100010001110000110010;
#10000;
data_in <= 24'b000111010010100000111110;
#10000;
data_in <= 24'b001011110011101001001110;
#10000;
data_in <= 24'b001110010100010001011000;
#10000;
data_in <= 24'b001101000100000001010010;
#10000;
data_in <= 24'b001010000011010001000110;
#10000;
data_in <= 24'b000111100010110000111110;
#10000;
data_in <= 24'b000100010001101000101110;
#10000;
data_in <= 24'b000100110001110000110000;
#10000;
data_in <= 24'b000110110010010000111000;
#10000;
data_in <= 24'b001001010010111101000001;
#10000;
data_in <= 24'b001010100011010001000110;
#10000;
data_in <= 24'b001001100011000001000001;
#10000;
data_in <= 24'b000111100010100000111001;
#10000;
data_in <= 24'b000110000010010100110101;
#10000;
data_in <= 24'b000110000001111100110010;
#10000;
data_in <= 24'b000110000001111100110010;
#10000;
data_in <= 24'b000110100010000100110100;
#10000;
data_in <= 24'b000111100010011000110111;
#10000;
data_in <= 24'b000111110010011100111000;
#10000;
data_in <= 24'b000110100010001100110001;
#10000;
data_in <= 24'b000101010001111000101100;
#10000;
data_in <= 24'b000100000001101000101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010100010110011010000010;
#10000;
data_in <= 24'b010101010110011110000100;
#10000;
data_in <= 24'b010110000110110010001011;
#10000;
data_in <= 24'b010000010101010001110101;
#10000;
data_in <= 24'b000011110010001001000101;
#10000;
data_in <= 24'b000000000001001100111000;
#10000;
data_in <= 24'b001001010011100001011110;
#10000;
data_in <= 24'b010010010101110110000110;
#10000;
data_in <= 24'b010000100101010001110001;
#10000;
data_in <= 24'b010110000110101010001001;
#10000;
data_in <= 24'b010111110111000110010000;
#10000;
data_in <= 24'b010011100110000110000010;
#10000;
data_in <= 24'b001101000100100001101011;
#10000;
data_in <= 24'b000111000010111101010100;
#10000;
data_in <= 24'b001000110011100001011110;
#10000;
data_in <= 24'b010001100101101010000011;
#10000;
data_in <= 24'b001010100011110101011000;
#10000;
data_in <= 24'b010011100110000001111101;
#10000;
data_in <= 24'b010101100110100010000111;
#10000;
data_in <= 24'b010100010110010010000101;
#10000;
data_in <= 24'b010100110110100010001000;
#10000;
data_in <= 24'b001110010100110101110000;
#10000;
data_in <= 24'b001010100100000001100100;
#10000;
data_in <= 24'b010001100101101110000001;
#10000;
data_in <= 24'b000110110010110001000110;
#10000;
data_in <= 24'b001101100100011101100010;
#10000;
data_in <= 24'b001111110101000101101110;
#10000;
data_in <= 24'b010001110101100101111000;
#10000;
data_in <= 24'b010100010110010110000100;
#10000;
data_in <= 24'b010001010101101001111010;
#10000;
data_in <= 24'b001110100100111001110001;
#10000;
data_in <= 24'b010001100101110001111111;
#10000;
data_in <= 24'b000101110010011100111110;
#10000;
data_in <= 24'b000111100010111101001001;
#10000;
data_in <= 24'b001011110100001101011100;
#10000;
data_in <= 24'b001111000100111101101010;
#10000;
data_in <= 24'b001111110101010001110000;
#10000;
data_in <= 24'b010000110101100001110111;
#10000;
data_in <= 24'b010001000101100101111000;
#10000;
data_in <= 24'b001111110101010001110100;
#10000;
data_in <= 24'b000101110010100000111101;
#10000;
data_in <= 24'b000110100010110001000011;
#10000;
data_in <= 24'b001011110100000101011000;
#10000;
data_in <= 24'b001110100100111001100111;
#10000;
data_in <= 24'b001101110100101001100101;
#10000;
data_in <= 24'b001111100101001101101111;
#10000;
data_in <= 24'b010000110101100001110100;
#10000;
data_in <= 24'b001100110100100101100101;
#10000;
data_in <= 24'b000101000010001100110110;
#10000;
data_in <= 24'b001000110011011001001011;
#10000;
data_in <= 24'b001100010100010001011001;
#10000;
data_in <= 24'b001100100100011101011101;
#10000;
data_in <= 24'b001101100100101001100011;
#10000;
data_in <= 24'b001110000100110101101000;
#10000;
data_in <= 24'b001101010100101001100101;
#10000;
data_in <= 24'b001100100100011101100010;
#10000;
data_in <= 24'b000011010001110100101110;
#10000;
data_in <= 24'b001011100011111101010010;
#10000;
data_in <= 24'b001011110100001001010111;
#10000;
data_in <= 24'b001010000011101101010000;
#10000;
data_in <= 24'b001110000100101001100001;
#10000;
data_in <= 24'b001101010100101001100000;
#10000;
data_in <= 24'b001011000100000001011001;
#10000;
data_in <= 24'b001110000100110101100011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b010000110101011110000000;
#10000;
data_in <= 24'b010000000101001101111110;
#10000;
data_in <= 24'b001111010101000001111011;
#10000;
data_in <= 24'b001110100100111001110111;
#10000;
data_in <= 24'b010011110110001110001100;
#10000;
data_in <= 24'b010111100111000010011001;
#10000;
data_in <= 24'b010110010110101110010100;
#10000;
data_in <= 24'b011001100111110010100101;
#10000;
data_in <= 24'b010010100110000010001001;
#10000;
data_in <= 24'b010010100110000010001001;
#10000;
data_in <= 24'b010010110101111010001001;
#10000;
data_in <= 24'b001110110100111101111000;
#10000;
data_in <= 24'b010000010101001101111100;
#10000;
data_in <= 24'b010100100110010110001011;
#10000;
data_in <= 24'b010110010110101010010001;
#10000;
data_in <= 24'b011001100111101010100011;
#10000;
data_in <= 24'b010110010110111010010100;
#10000;
data_in <= 24'b011000010111011010011100;
#10000;
data_in <= 24'b011010100111110010100101;
#10000;
data_in <= 24'b010011000101111110000101;
#10000;
data_in <= 24'b001110000100100101110000;
#10000;
data_in <= 24'b010001110101100101111110;
#10000;
data_in <= 24'b010110000110100010001101;
#10000;
data_in <= 24'b010111110111001010011000;
#10000;
data_in <= 24'b010110110111000110010101;
#10000;
data_in <= 24'b011011001000001010100110;
#10000;
data_in <= 24'b100000011001010010111001;
#10000;
data_in <= 24'b010111110111001010010111;
#10000;
data_in <= 24'b001110010100110001101111;
#10000;
data_in <= 24'b010000110101011001111001;
#10000;
data_in <= 24'b010101010110011010000111;
#10000;
data_in <= 24'b010101100110101010001101;
#10000;
data_in <= 24'b010010110101111110000010;
#10000;
data_in <= 24'b010111000111000010010011;
#10000;
data_in <= 24'b011100111000011010100111;
#10000;
data_in <= 24'b010101100110100110001010;
#10000;
data_in <= 24'b001100110100010101100100;
#10000;
data_in <= 24'b001111010100111101101110;
#10000;
data_in <= 24'b010100010110000101111110;
#10000;
data_in <= 24'b010101010110100110001000;
#10000;
data_in <= 24'b001101010100101001101001;
#10000;
data_in <= 24'b001110010100110101101100;
#10000;
data_in <= 24'b010001000101100101110101;
#10000;
data_in <= 24'b001100010100001101100000;
#10000;
data_in <= 24'b000111010011000001001011;
#10000;
data_in <= 24'b001010010011101001010101;
#10000;
data_in <= 24'b001110110100110001100110;
#10000;
data_in <= 24'b010011110110001001111101;
#10000;
data_in <= 24'b001011010100001001011101;
#10000;
data_in <= 24'b001000010011010001001111;
#10000;
data_in <= 24'b000110010010110101000110;
#10000;
data_in <= 24'b000011010001111000111000;
#10000;
data_in <= 24'b000001110001100100110000;
#10000;
data_in <= 24'b000010110001101100110010;
#10000;
data_in <= 24'b000101010010011000111011;
#10000;
data_in <= 24'b001101100100011001011101;
#10000;
data_in <= 24'b001101000100100001100001;
#10000;
data_in <= 24'b000111000010111001000101;
#10000;
data_in <= 24'b000001110001100100110000;
#10000;
data_in <= 24'b000000000000111100100100;
#10000;
data_in <= 24'b000000000001000000100011;
#10000;
data_in <= 24'b000000000000011000011001;
#10000;
data_in <= 24'b000000000000001100010101;
#10000;
data_in <= 24'b000110000010011100111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011001011000001110101100;
#10000;
data_in <= 24'b011001001000011010110001;
#10000;
data_in <= 24'b011010101000101010110101;
#10000;
data_in <= 24'b011010101000110010110111;
#10000;
data_in <= 24'b011010101000110010110111;
#10000;
data_in <= 24'b011010111000111010110110;
#10000;
data_in <= 24'b011011101001000110111001;
#10000;
data_in <= 24'b011100101001010110111101;
#10000;
data_in <= 24'b011000000111110010100101;
#10000;
data_in <= 24'b010111010111111110101010;
#10000;
data_in <= 24'b011001011000010110110000;
#10000;
data_in <= 24'b011001111000100110110100;
#10000;
data_in <= 24'b011010011000110010110100;
#10000;
data_in <= 24'b011010101000110110110101;
#10000;
data_in <= 24'b011010111000111110110101;
#10000;
data_in <= 24'b011011011001000110110111;
#10000;
data_in <= 24'b010111010111011110011111;
#10000;
data_in <= 24'b010110110111101110100100;
#10000;
data_in <= 24'b011001001000001010101011;
#10000;
data_in <= 24'b011001111000011110110000;
#10000;
data_in <= 24'b011010111000101110110100;
#10000;
data_in <= 24'b011011011000110110110110;
#10000;
data_in <= 24'b011011011000110110110110;
#10000;
data_in <= 24'b011011001000110110110100;
#10000;
data_in <= 24'b010110110111010110011010;
#10000;
data_in <= 24'b010111000111100110100000;
#10000;
data_in <= 24'b011000010111111010100101;
#10000;
data_in <= 24'b011001001000001110101010;
#10000;
data_in <= 24'b011010011000011110110000;
#10000;
data_in <= 24'b011011011000101110110100;
#10000;
data_in <= 24'b011011011000101110110100;
#10000;
data_in <= 24'b011010001000100010110001;
#10000;
data_in <= 24'b010110000111000010010100;
#10000;
data_in <= 24'b010110100111010110011010;
#10000;
data_in <= 24'b010111100111100110011110;
#10000;
data_in <= 24'b010111110111101010011111;
#10000;
data_in <= 24'b011000110111110110100101;
#10000;
data_in <= 24'b011010001000010110101100;
#10000;
data_in <= 24'b011010101000011110101110;
#10000;
data_in <= 24'b011001101000010110101100;
#10000;
data_in <= 24'b010101100110101110001011;
#10000;
data_in <= 24'b010110110111010010010110;
#10000;
data_in <= 24'b011000000111100010011100;
#10000;
data_in <= 24'b010111110111011110011011;
#10000;
data_in <= 24'b010111110111100110011101;
#10000;
data_in <= 24'b011001101000000110100110;
#10000;
data_in <= 24'b011011001000011110101100;
#10000;
data_in <= 24'b011010011000011010101101;
#10000;
data_in <= 24'b010011000101111001111011;
#10000;
data_in <= 24'b010110000110110010001011;
#10000;
data_in <= 24'b011000000111010110010101;
#10000;
data_in <= 24'b010111110111010010010100;
#10000;
data_in <= 24'b010111110111010110011000;
#10000;
data_in <= 24'b011001010111110110100001;
#10000;
data_in <= 24'b011010101000010010101001;
#10000;
data_in <= 24'b011010101000010010101100;
#10000;
data_in <= 24'b001111110100111001101000;
#10000;
data_in <= 24'b010011110110000001111011;
#10000;
data_in <= 24'b010110100110110010001001;
#10000;
data_in <= 24'b010110010110111010001010;
#10000;
data_in <= 24'b010110010110110110001100;
#10000;
data_in <= 24'b010111100111010110010101;
#10000;
data_in <= 24'b011001100111110010011111;
#10000;
data_in <= 24'b011000110111110110100010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011101101001011010111111;
#10000;
data_in <= 24'b011101111001100010111111;
#10000;
data_in <= 24'b011110001001100111000000;
#10000;
data_in <= 24'b011110101001101111000010;
#10000;
data_in <= 24'b011110111001110011000011;
#10000;
data_in <= 24'b011110111001110011000011;
#10000;
data_in <= 24'b011111001001111011000010;
#10000;
data_in <= 24'b011111001001110111000100;
#10000;
data_in <= 24'b011101011001011010111101;
#10000;
data_in <= 24'b011101011001011110111011;
#10000;
data_in <= 24'b011101101001100010111100;
#10000;
data_in <= 24'b011110001001101110111101;
#10000;
data_in <= 24'b011110001001101010111110;
#10000;
data_in <= 24'b011110011001110010111110;
#10000;
data_in <= 24'b011110011001110010111110;
#10000;
data_in <= 24'b011110011001110010111110;
#10000;
data_in <= 24'b011100101001001110111010;
#10000;
data_in <= 24'b011100101001001110111010;
#10000;
data_in <= 24'b011100011001010110111011;
#10000;
data_in <= 24'b011100101001011010111010;
#10000;
data_in <= 24'b011100101001011010111100;
#10000;
data_in <= 24'b011100111001011110111011;
#10000;
data_in <= 24'b011100111001011110111011;
#10000;
data_in <= 24'b011100111001011110111011;
#10000;
data_in <= 24'b011011101000111110110110;
#10000;
data_in <= 24'b011011101000111110110110;
#10000;
data_in <= 24'b011011001001000010110110;
#10000;
data_in <= 24'b011011011001000010111000;
#10000;
data_in <= 24'b011011011001000010111000;
#10000;
data_in <= 24'b011011101001000110111001;
#10000;
data_in <= 24'b011011111001001010111010;
#10000;
data_in <= 24'b011011111001001010111010;
#10000;
data_in <= 24'b011010101000101010110011;
#10000;
data_in <= 24'b011010101000101010110011;
#10000;
data_in <= 24'b011010001000101110110011;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011010001000101110110110;
#10000;
data_in <= 24'b011010011000110010110111;
#10000;
data_in <= 24'b011010101000110110111000;
#10000;
data_in <= 24'b011010111000111010111001;
#10000;
data_in <= 24'b011010001000011010101111;
#10000;
data_in <= 24'b011001101000011010101111;
#10000;
data_in <= 24'b011001101000011010110001;
#10000;
data_in <= 24'b011001001000011010110001;
#10000;
data_in <= 24'b011001001000011110110011;
#10000;
data_in <= 24'b011001101000100110110101;
#10000;
data_in <= 24'b011001101000101110110111;
#10000;
data_in <= 24'b011010011000110010111000;
#10000;
data_in <= 24'b011001111000001110101100;
#10000;
data_in <= 24'b011001011000001110101100;
#10000;
data_in <= 24'b011000111000001110101110;
#10000;
data_in <= 24'b011000011000001010101111;
#10000;
data_in <= 24'b011000101000010010110010;
#10000;
data_in <= 24'b011001011000011110110101;
#10000;
data_in <= 24'b011001111000100110110111;
#10000;
data_in <= 24'b011010011000110010111000;
#10000;
data_in <= 24'b011010001000001010101010;
#10000;
data_in <= 24'b011001011000000110101010;
#10000;
data_in <= 24'b011000111000000010101100;
#10000;
data_in <= 24'b011000101000000110101110;
#10000;
data_in <= 24'b011000101000001110110000;
#10000;
data_in <= 24'b011001011000011010110100;
#10000;
data_in <= 24'b011010001000100110110111;
#10000;
data_in <= 24'b011010101000101110111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011011101000111010111001;
#10000;
data_in <= 24'b011000011000000010101101;
#10000;
data_in <= 24'b010100110111000110100000;
#10000;
data_in <= 24'b010010100110101010011011;
#10000;
data_in <= 24'b010010010110100010011011;
#10000;
data_in <= 24'b010011000110101110100000;
#10000;
data_in <= 24'b010100110111001010100111;
#10000;
data_in <= 24'b010110100111100110101110;
#10000;
data_in <= 24'b011101101001011110111110;
#10000;
data_in <= 24'b011010111000111010110110;
#10000;
data_in <= 24'b011000101000010010101111;
#10000;
data_in <= 24'b011000001000001110101111;
#10000;
data_in <= 24'b011000101000010010110010;
#10000;
data_in <= 24'b011001011000011010110111;
#10000;
data_in <= 24'b011010111000110010111101;
#10000;
data_in <= 24'b011100011001001011000011;
#10000;
data_in <= 24'b011101001001100010111110;
#10000;
data_in <= 24'b011100001001001110111011;
#10000;
data_in <= 24'b011011101001000010111011;
#10000;
data_in <= 24'b011100001001001110111111;
#10000;
data_in <= 24'b011101001001011011000100;
#10000;
data_in <= 24'b011101011001100111000111;
#10000;
data_in <= 24'b011110101001111011001110;
#10000;
data_in <= 24'b011111101010001011010010;
#10000;
data_in <= 24'b011100001001010010111010;
#10000;
data_in <= 24'b011011101001001010111000;
#10000;
data_in <= 24'b011011101001001010111010;
#10000;
data_in <= 24'b011101001001011111000010;
#10000;
data_in <= 24'b011101111001110011001000;
#10000;
data_in <= 24'b011110011001110111001011;
#10000;
data_in <= 24'b011111101010001011010010;
#10000;
data_in <= 24'b100000101010011011010100;
#10000;
data_in <= 24'b011100001001001110111011;
#10000;
data_in <= 24'b011011111001001110111001;
#10000;
data_in <= 24'b011100001001010010111100;
#10000;
data_in <= 24'b011101101001100111000100;
#10000;
data_in <= 24'b011110011001111011001010;
#10000;
data_in <= 24'b011111011010001011001110;
#10000;
data_in <= 24'b100000101010100111010110;
#10000;
data_in <= 24'b100010001010111111011100;
#10000;
data_in <= 24'b011011111001001010111010;
#10000;
data_in <= 24'b011011101001001010111000;
#10000;
data_in <= 24'b011100001001010010111100;
#10000;
data_in <= 24'b011101101001101011000010;
#10000;
data_in <= 24'b011110101010000011001010;
#10000;
data_in <= 24'b011111111010010011010000;
#10000;
data_in <= 24'b100001011010110011011001;
#10000;
data_in <= 24'b100011011011010011100001;
#10000;
data_in <= 24'b011011001000111110110111;
#10000;
data_in <= 24'b011011001001000010110110;
#10000;
data_in <= 24'b011011111001001110111011;
#10000;
data_in <= 24'b011101001001100011000000;
#10000;
data_in <= 24'b011101101001110011000110;
#10000;
data_in <= 24'b011110101010000011001010;
#10000;
data_in <= 24'b011111111010011011010010;
#10000;
data_in <= 24'b100001111010111011011010;
#10000;
data_in <= 24'b011011101001001010111000;
#10000;
data_in <= 24'b011011101001001010110110;
#10000;
data_in <= 24'b011100011001010110111011;
#10000;
data_in <= 24'b011101011001100111000001;
#10000;
data_in <= 24'b011101101001100111000100;
#10000;
data_in <= 24'b011101011001101111000101;
#10000;
data_in <= 24'b011110001001111111001011;
#10000;
data_in <= 24'b011111111010011011010010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011010101000011110111010;
#10000;
data_in <= 24'b011101111001010111000100;
#10000;
data_in <= 24'b100010011010011011010010;
#10000;
data_in <= 24'b100101111011011011011101;
#10000;
data_in <= 24'b101001101100010011100111;
#10000;
data_in <= 24'b101100011101000011101111;
#10000;
data_in <= 24'b101101101101011111110001;
#10000;
data_in <= 24'b101101101101100011110000;
#10000;
data_in <= 24'b011110011001101011001000;
#10000;
data_in <= 24'b100001001010010111010010;
#10000;
data_in <= 24'b100101001011010011011101;
#10000;
data_in <= 24'b100111111100000111100101;
#10000;
data_in <= 24'b101010111100110011101101;
#10000;
data_in <= 24'b101101111101011111110100;
#10000;
data_in <= 24'b101111101101110011110111;
#10000;
data_in <= 24'b101111011101110111110100;
#10000;
data_in <= 24'b100010011010101111011001;
#10000;
data_in <= 24'b100100101011010111100001;
#10000;
data_in <= 24'b100111101100000111101001;
#10000;
data_in <= 24'b101001111100100111101101;
#10000;
data_in <= 24'b101100001101000011110011;
#10000;
data_in <= 24'b101110001101101011111000;
#10000;
data_in <= 24'b101111011101110111111010;
#10000;
data_in <= 24'b101111101101110111110110;
#10000;
data_in <= 24'b100100011011001111100001;
#10000;
data_in <= 24'b100110001011101111100111;
#10000;
data_in <= 24'b101000011100010011101100;
#10000;
data_in <= 24'b101001011100100111101101;
#10000;
data_in <= 24'b101011001100111111110001;
#10000;
data_in <= 24'b101101001101010111110110;
#10000;
data_in <= 24'b101110011101100111110110;
#10000;
data_in <= 24'b101110001101100111110011;
#10000;
data_in <= 24'b100100001011010011100010;
#10000;
data_in <= 24'b100101111011110011101000;
#10000;
data_in <= 24'b100111111100001111101011;
#10000;
data_in <= 24'b101000111100011111101101;
#10000;
data_in <= 24'b101010011100101111101111;
#10000;
data_in <= 24'b101011111101001011110011;
#10000;
data_in <= 24'b101100111101010111110011;
#10000;
data_in <= 24'b101100111101010111110010;
#10000;
data_in <= 24'b100011111011010011100000;
#10000;
data_in <= 24'b100101101011110011100110;
#10000;
data_in <= 24'b100111111100001011101101;
#10000;
data_in <= 24'b101000101100011111101101;
#10000;
data_in <= 24'b101001111100101111101111;
#10000;
data_in <= 24'b101011101101000111110011;
#10000;
data_in <= 24'b101100101101001111110100;
#10000;
data_in <= 24'b101100011101001111110001;
#10000;
data_in <= 24'b100010101011000111011101;
#10000;
data_in <= 24'b100100011011100111100011;
#10000;
data_in <= 24'b100110101100000011101010;
#10000;
data_in <= 24'b100111111100010011101010;
#10000;
data_in <= 24'b101001001100100011101100;
#10000;
data_in <= 24'b101010001100110111101111;
#10000;
data_in <= 24'b101011001100111111110001;
#10000;
data_in <= 24'b101010101100110111101111;
#10000;
data_in <= 24'b100001011010110011011000;
#10000;
data_in <= 24'b100011001011010011011110;
#10000;
data_in <= 24'b100101101011110011100110;
#10000;
data_in <= 24'b100110011100000011100111;
#10000;
data_in <= 24'b100111101100001111101001;
#10000;
data_in <= 24'b101000111100011111101011;
#10000;
data_in <= 24'b101001101100100011101100;
#10000;
data_in <= 24'b101001001100011011101010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b101111001101110111110001;
#10000;
data_in <= 24'b101111001101110111110001;
#10000;
data_in <= 24'b101110011101101111110011;
#10000;
data_in <= 24'b101101111101100111110110;
#10000;
data_in <= 24'b101100011101011011111000;
#10000;
data_in <= 24'b101001111100110011110010;
#10000;
data_in <= 24'b100110101100000011101010;
#10000;
data_in <= 24'b100011111011011011100011;
#10000;
data_in <= 24'b101111101101110111110010;
#10000;
data_in <= 24'b101111111101111011110011;
#10000;
data_in <= 24'b101111111101111011110111;
#10000;
data_in <= 24'b101111011101110111111010;
#10000;
data_in <= 24'b101101001101011111111001;
#10000;
data_in <= 24'b101001101100101111110001;
#10000;
data_in <= 24'b100101111011110011101000;
#10000;
data_in <= 24'b100011001011001111100000;
#10000;
data_in <= 24'b101111011101110011110011;
#10000;
data_in <= 24'b110000001101111111110110;
#10000;
data_in <= 24'b110000011101111111111010;
#10000;
data_in <= 24'b101110111101110111111011;
#10000;
data_in <= 24'b101100011101010011110110;
#10000;
data_in <= 24'b101000011100010111101101;
#10000;
data_in <= 24'b100100101011011111100011;
#10000;
data_in <= 24'b100001111010111011011011;
#10000;
data_in <= 24'b101110101101100111110010;
#10000;
data_in <= 24'b101111001101101111110100;
#10000;
data_in <= 24'b101110111101101111111000;
#10000;
data_in <= 24'b101101011101011011110111;
#10000;
data_in <= 24'b101010001100110011110000;
#10000;
data_in <= 24'b100110111011111111100111;
#10000;
data_in <= 24'b100011011011001011011110;
#10000;
data_in <= 24'b100001001010101111011000;
#10000;
data_in <= 24'b101101111101011111110100;
#10000;
data_in <= 24'b101101001101011011110011;
#10000;
data_in <= 24'b101100011101001011110011;
#10000;
data_in <= 24'b101010101100110111101111;
#10000;
data_in <= 24'b100111111100001111101001;
#10000;
data_in <= 24'b100101001011011111100010;
#10000;
data_in <= 24'b100010001010110111011001;
#10000;
data_in <= 24'b100000101010011011010100;
#10000;
data_in <= 24'b101100011101001111110001;
#10000;
data_in <= 24'b101010111100111011101111;
#10000;
data_in <= 24'b101001001100011111101001;
#10000;
data_in <= 24'b100111001100000011100110;
#10000;
data_in <= 24'b100101001011100011100000;
#10000;
data_in <= 24'b100010111010111011011010;
#10000;
data_in <= 24'b100000011010001111010001;
#10000;
data_in <= 24'b011110101001110011001010;
#10000;
data_in <= 24'b101001101100100111101011;
#10000;
data_in <= 24'b100111011100000111100101;
#10000;
data_in <= 24'b100101011011100111011111;
#10000;
data_in <= 24'b100011111011001011011010;
#10000;
data_in <= 24'b100010011010110011010111;
#10000;
data_in <= 24'b011111111010001011001110;
#10000;
data_in <= 24'b011100011001001111000001;
#10000;
data_in <= 24'b011010001000100110110111;
#10000;
data_in <= 24'b100110111011111111100011;
#10000;
data_in <= 24'b100100111011011111011101;
#10000;
data_in <= 24'b100010101010110111010101;
#10000;
data_in <= 24'b100001011010011111010010;
#10000;
data_in <= 24'b100000001010001111001111;
#10000;
data_in <= 24'b011101011001100011000100;
#10000;
data_in <= 24'b011001011000011010110100;
#10000;
data_in <= 24'b010110010111011110100110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100001011010110111011101;
#10000;
data_in <= 24'b100000101010100011011000;
#10000;
data_in <= 24'b011111001010000011001110;
#10000;
data_in <= 24'b011101101001100111000101;
#10000;
data_in <= 24'b011100111001010111000000;
#10000;
data_in <= 24'b011011001000110010110101;
#10000;
data_in <= 24'b010110010111100010011111;
#10000;
data_in <= 24'b010010100110011010001001;
#10000;
data_in <= 24'b100000111010101111011100;
#10000;
data_in <= 24'b011111111010010011010110;
#10000;
data_in <= 24'b011110011001110111001101;
#10000;
data_in <= 24'b011101001001011011000100;
#10000;
data_in <= 24'b011100101001001010111101;
#10000;
data_in <= 24'b011001111000010110101110;
#10000;
data_in <= 24'b010011110110110010010001;
#10000;
data_in <= 24'b001110100101010101110111;
#10000;
data_in <= 24'b100000101010011111011001;
#10000;
data_in <= 24'b011111011010001011010100;
#10000;
data_in <= 24'b011110001001110011001100;
#10000;
data_in <= 24'b011100111001011011000010;
#10000;
data_in <= 24'b011011111000111110111000;
#10000;
data_in <= 24'b010111110111111010100101;
#10000;
data_in <= 24'b010000110110000010000101;
#10000;
data_in <= 24'b001011110100100001101010;
#10000;
data_in <= 24'b011110111010000111010001;
#10000;
data_in <= 24'b011110011001110111001101;
#10000;
data_in <= 24'b011101001001011011000100;
#10000;
data_in <= 24'b011011011000111110111010;
#10000;
data_in <= 24'b011001001000001010101011;
#10000;
data_in <= 24'b010100010110111010010011;
#10000;
data_in <= 24'b001110010101010101111000;
#10000;
data_in <= 24'b001010100100000101100001;
#10000;
data_in <= 24'b011100111001011111000101;
#10000;
data_in <= 24'b011100001001001011000000;
#10000;
data_in <= 24'b011010111000101010110111;
#10000;
data_in <= 24'b011000010111111110101000;
#10000;
data_in <= 24'b010100110110110110010101;
#10000;
data_in <= 24'b001111100101100001111100;
#10000;
data_in <= 24'b001011000100010101100101;
#10000;
data_in <= 24'b001001000011100101011000;
#10000;
data_in <= 24'b011011001000111010111100;
#10000;
data_in <= 24'b011001011000011010110011;
#10000;
data_in <= 24'b010111010111101010100110;
#10000;
data_in <= 24'b010100000110110110010100;
#10000;
data_in <= 24'b010000010101101110000000;
#10000;
data_in <= 24'b001011110100100001101010;
#10000;
data_in <= 24'b001000100011101001011000;
#10000;
data_in <= 24'b000111100011001101001111;
#10000;
data_in <= 24'b010111000111110110101010;
#10000;
data_in <= 24'b010100000110111110011100;
#10000;
data_in <= 24'b010001000110000010001001;
#10000;
data_in <= 24'b001110110101011001111011;
#10000;
data_in <= 24'b001100100100101001101110;
#10000;
data_in <= 24'b001001100011110101011101;
#10000;
data_in <= 24'b000110110011000101001101;
#10000;
data_in <= 24'b000110000010101101000110;
#10000;
data_in <= 24'b010010000110011110010100;
#10000;
data_in <= 24'b001110000101010110000001;
#10000;
data_in <= 24'b001010100100001101101101;
#10000;
data_in <= 24'b001001010011111101100100;
#10000;
data_in <= 24'b001001100011110001011111;
#10000;
data_in <= 24'b000111110011010001010011;
#10000;
data_in <= 24'b000100110010100001000100;
#10000;
data_in <= 24'b000011010010000100111010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101100100111001101100;
#10000;
data_in <= 24'b001011110100010001100000;
#10000;
data_in <= 24'b001000100011010101010000;
#10000;
data_in <= 24'b000101110010100001000010;
#10000;
data_in <= 24'b000100110010000100111000;
#10000;
data_in <= 24'b000011110001110100110000;
#10000;
data_in <= 24'b000011100001100000101010;
#10000;
data_in <= 24'b000011000001010000100101;
#10000;
data_in <= 24'b001100110100011101100110;
#10000;
data_in <= 24'b001011000011110101011000;
#10000;
data_in <= 24'b000111100010110101000111;
#10000;
data_in <= 24'b000101010010001100111010;
#10000;
data_in <= 24'b000100010001111000110100;
#10000;
data_in <= 24'b000100000001101100101111;
#10000;
data_in <= 24'b000011010001011100101001;
#10000;
data_in <= 24'b000010110001010000100010;
#10000;
data_in <= 24'b001010110011110101011100;
#10000;
data_in <= 24'b001000110011000101001101;
#10000;
data_in <= 24'b000101000010001100111101;
#10000;
data_in <= 24'b000011100001110000110011;
#10000;
data_in <= 24'b000011010001101000110000;
#10000;
data_in <= 24'b000011110001101100101101;
#10000;
data_in <= 24'b000011010001011100101000;
#10000;
data_in <= 24'b000010110001010000100010;
#10000;
data_in <= 24'b001000010011001101010000;
#10000;
data_in <= 24'b000110010010100001000010;
#10000;
data_in <= 24'b000011100001110000110011;
#10000;
data_in <= 24'b000010010001011000101100;
#10000;
data_in <= 24'b000011010001100000101100;
#10000;
data_in <= 24'b000100010001101100101101;
#10000;
data_in <= 24'b000100000001100000101001;
#10000;
data_in <= 24'b000011000001010100100010;
#10000;
data_in <= 24'b000110010010101001000101;
#10000;
data_in <= 24'b000101000010001000111001;
#10000;
data_in <= 24'b000010110001011100101111;
#10000;
data_in <= 24'b000010000001010100101011;
#10000;
data_in <= 24'b000011010001100000101100;
#10000;
data_in <= 24'b000100100001110000101101;
#10000;
data_in <= 24'b000100110001110000101010;
#10000;
data_in <= 24'b000100000001100100100110;
#10000;
data_in <= 24'b000100110010001000111100;
#10000;
data_in <= 24'b000011110001110100110011;
#10000;
data_in <= 24'b000010110001100000101110;
#10000;
data_in <= 24'b000010110001011000101010;
#10000;
data_in <= 24'b000100000001101000101100;
#10000;
data_in <= 24'b000100100001110000101101;
#10000;
data_in <= 24'b000101000001110100101011;
#10000;
data_in <= 24'b000100110001110000101001;
#10000;
data_in <= 24'b000011000001110000110011;
#10000;
data_in <= 24'b000011100001101100110001;
#10000;
data_in <= 24'b000011100001100100101111;
#10000;
data_in <= 24'b000011010001100000101100;
#10000;
data_in <= 24'b000100000001101000101100;
#10000;
data_in <= 24'b000100010001101100101100;
#10000;
data_in <= 24'b000100100001110100101011;
#10000;
data_in <= 24'b000100110001111100101011;
#10000;
data_in <= 24'b000010100001100000101111;
#10000;
data_in <= 24'b000011000001100100101111;
#10000;
data_in <= 24'b000011110001101000101110;
#10000;
data_in <= 24'b000011110001101100101101;
#10000;
data_in <= 24'b000100000001101000101100;
#10000;
data_in <= 24'b000100000001101100101001;
#10000;
data_in <= 24'b000100100001110100101011;
#10000;
data_in <= 24'b000100110001111100101011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000011100001010100100100;
#10000;
data_in <= 24'b000100010001100000100111;
#10000;
data_in <= 24'b000100110001100100100110;
#10000;
data_in <= 24'b000100100001100000100101;
#10000;
data_in <= 24'b000101010001101100101000;
#10000;
data_in <= 24'b000110010001111100101100;
#10000;
data_in <= 24'b000101100001111000101011;
#10000;
data_in <= 24'b000100100001101000100111;
#10000;
data_in <= 24'b000011010001010000100011;
#10000;
data_in <= 24'b000100010001100100100110;
#10000;
data_in <= 24'b000100100001101000100111;
#10000;
data_in <= 24'b000100010001100100100110;
#10000;
data_in <= 24'b000100110001101100101000;
#10000;
data_in <= 24'b000101110010000000101101;
#10000;
data_in <= 24'b000110010010001000101111;
#10000;
data_in <= 24'b000110000010000100101110;
#10000;
data_in <= 24'b000011000001010100100011;
#10000;
data_in <= 24'b000100000001100100100110;
#10000;
data_in <= 24'b000100110001110000101001;
#10000;
data_in <= 24'b000100100001110000100110;
#10000;
data_in <= 24'b000100110001110000101001;
#10000;
data_in <= 24'b000110000010000100101110;
#10000;
data_in <= 24'b000111010010011000110011;
#10000;
data_in <= 24'b000111100010101000110110;
#10000;
data_in <= 24'b000011010001011000100011;
#10000;
data_in <= 24'b000100010001101000100111;
#10000;
data_in <= 24'b000100110001110100100111;
#10000;
data_in <= 24'b000100100001110000100110;
#10000;
data_in <= 24'b000100100001101100101000;
#10000;
data_in <= 24'b000101000010000000101100;
#10000;
data_in <= 24'b000110110010011100110011;
#10000;
data_in <= 24'b000111110010110100111001;
#10000;
data_in <= 24'b000100010001101000100111;
#10000;
data_in <= 24'b000100100001110000100110;
#10000;
data_in <= 24'b000100010001110100100111;
#10000;
data_in <= 24'b000100000001110000100110;
#10000;
data_in <= 24'b000011110001101100100101;
#10000;
data_in <= 24'b000011100001110100100110;
#10000;
data_in <= 24'b000101010010010000101101;
#10000;
data_in <= 24'b000110100010101100110100;
#10000;
data_in <= 24'b000101000001111000101000;
#10000;
data_in <= 24'b000100010001110100100111;
#10000;
data_in <= 24'b000100000001110000100110;
#10000;
data_in <= 24'b000011100001110100100110;
#10000;
data_in <= 24'b000011010001110000100101;
#10000;
data_in <= 24'b000010110001110000100101;
#10000;
data_in <= 24'b000100000010000100101010;
#10000;
data_in <= 24'b000101010010100000110000;
#10000;
data_in <= 24'b000101010010000100101011;
#10000;
data_in <= 24'b000100010001110100100111;
#10000;
data_in <= 24'b000011110001110000100100;
#10000;
data_in <= 24'b000011110001111100100110;
#10000;
data_in <= 24'b000011010001111000100111;
#10000;
data_in <= 24'b000010110001111000100110;
#10000;
data_in <= 24'b000011010001111100101010;
#10000;
data_in <= 24'b000100000010010000101111;
#10000;
data_in <= 24'b000101110010001100101101;
#10000;
data_in <= 24'b000100010001110100100111;
#10000;
data_in <= 24'b000011000001110000100011;
#10000;
data_in <= 24'b000011100010000000100111;
#10000;
data_in <= 24'b000011100010000100101001;
#10000;
data_in <= 24'b000011010010000000101000;
#10000;
data_in <= 24'b000011000010000000101011;
#10000;
data_in <= 24'b000011110010001100101110;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000100100001101100100100;
#10000;
data_in <= 24'b000100010001101000100011;
#10000;
data_in <= 24'b000100110001110000100110;
#10000;
data_in <= 24'b000101000001110000101001;
#10000;
data_in <= 24'b000100000001011100100110;
#10000;
data_in <= 24'b000010100001000100100000;
#10000;
data_in <= 24'b000010110001001000100011;
#10000;
data_in <= 24'b000100010001100000101001;
#10000;
data_in <= 24'b000010100001010100011101;
#10000;
data_in <= 24'b000010110001010100011111;
#10000;
data_in <= 24'b000011110001100100100011;
#10000;
data_in <= 24'b000100110001110000101001;
#10000;
data_in <= 24'b000100000001100100100111;
#10000;
data_in <= 24'b000010100001001000100011;
#10000;
data_in <= 24'b000001100000111000011111;
#10000;
data_in <= 24'b000010000000111100100010;
#10000;
data_in <= 24'b000011100001101000100100;
#10000;
data_in <= 24'b000011110001101100100101;
#10000;
data_in <= 24'b000100110001111100101011;
#10000;
data_in <= 24'b000110010010010000110010;
#10000;
data_in <= 24'b000110000010001100110001;
#10000;
data_in <= 24'b000100000001101000101011;
#10000;
data_in <= 24'b000010000001001000100100;
#10000;
data_in <= 24'b000001000000110100100001;
#10000;
data_in <= 24'b000100100010001000101110;
#10000;
data_in <= 24'b000100110010001100101111;
#10000;
data_in <= 24'b000101100010011000110011;
#10000;
data_in <= 24'b000111000010101100111011;
#10000;
data_in <= 24'b000111110010111000111110;
#10000;
data_in <= 24'b000111000010101000111100;
#10000;
data_in <= 24'b000101000010001000110101;
#10000;
data_in <= 24'b000011100001101100110001;
#10000;
data_in <= 24'b000111000010110100111010;
#10000;
data_in <= 24'b000111000010110000111100;
#10000;
data_in <= 24'b000111010010110100111101;
#10000;
data_in <= 24'b001000100011001001000011;
#10000;
data_in <= 24'b001001110011011001001001;
#10000;
data_in <= 24'b001010010011011101001101;
#10000;
data_in <= 24'b001001000011001001001000;
#10000;
data_in <= 24'b000111100010110001000011;
#10000;
data_in <= 24'b001101110100101101011100;
#10000;
data_in <= 24'b001101110100101101011100;
#10000;
data_in <= 24'b001101010100100101011010;
#10000;
data_in <= 24'b001100110100011101011001;
#10000;
data_in <= 24'b001100110100011001011011;
#10000;
data_in <= 24'b001100000100001001011001;
#10000;
data_in <= 24'b001010000011101001010001;
#10000;
data_in <= 24'b000111110011000001001010;
#10000;
data_in <= 24'b010011010110001101110101;
#10000;
data_in <= 24'b010100010110011101111001;
#10000;
data_in <= 24'b010100110110100101111011;
#10000;
data_in <= 24'b010011110110010001111001;
#10000;
data_in <= 24'b010010010101111001110011;
#10000;
data_in <= 24'b010000000101010101101011;
#10000;
data_in <= 24'b001100100100011001011111;
#10000;
data_in <= 24'b001001000011011101010010;
#10000;
data_in <= 24'b010010000110000001110010;
#10000;
data_in <= 24'b010100100110101001111100;
#10000;
data_in <= 24'b010110110111001110000111;
#10000;
data_in <= 24'b010111010111010110001001;
#10000;
data_in <= 24'b010110100111000110000111;
#10000;
data_in <= 24'b010100000110011101111101;
#10000;
data_in <= 24'b010000000101010101110000;
#10000;
data_in <= 24'b001100010100011001100001;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000100000001011000101001;
#10000;
data_in <= 24'b000101110001110100110000;
#10000;
data_in <= 24'b000111000010001100110100;
#10000;
data_in <= 24'b000110010010000000110001;
#10000;
data_in <= 24'b000100010001100000101001;
#10000;
data_in <= 24'b000010110001001000100001;
#10000;
data_in <= 24'b000011000001001100100010;
#10000;
data_in <= 24'b000011010001100000100110;
#10000;
data_in <= 24'b000011100001010100101000;
#10000;
data_in <= 24'b000100100001100100101100;
#10000;
data_in <= 24'b000101000001101100101110;
#10000;
data_in <= 24'b000100010001100100101010;
#10000;
data_in <= 24'b000010110001001100100100;
#10000;
data_in <= 24'b000010100001001100100001;
#10000;
data_in <= 24'b000100000001100100100111;
#10000;
data_in <= 24'b000101000001111100101101;
#10000;
data_in <= 24'b000100000001100100101101;
#10000;
data_in <= 24'b000100010001101000101110;
#10000;
data_in <= 24'b000100010001101000101110;
#10000;
data_in <= 24'b000011100001100000101010;
#10000;
data_in <= 24'b000011000001011000101000;
#10000;
data_in <= 24'b000011100001100000101001;
#10000;
data_in <= 24'b000101100010000000110001;
#10000;
data_in <= 24'b000110100010011100110111;
#10000;
data_in <= 24'b000101010010001000111000;
#10000;
data_in <= 24'b000101100010001100111001;
#10000;
data_in <= 24'b000101110010010000111010;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
data_in <= 24'b000101100010010000110111;
#10000;
data_in <= 24'b000101010010001100110101;
#10000;
data_in <= 24'b000101100010010000110110;
#10000;
data_in <= 24'b000101110010010100110111;
#10000;
data_in <= 24'b000110110010100101000000;
#10000;
data_in <= 24'b000111100010110001000011;
#10000;
data_in <= 24'b001000100011000001000111;
#10000;
data_in <= 24'b001001010011001101001001;
#10000;
data_in <= 24'b001001000011001001001000;
#10000;
data_in <= 24'b000111100010110101000000;
#10000;
data_in <= 24'b000101100010010100111000;
#10000;
data_in <= 24'b000011110001111000110001;
#10000;
data_in <= 24'b000111000010110101000111;
#10000;
data_in <= 24'b000111010010111001001000;
#10000;
data_in <= 24'b001000010011001001001100;
#10000;
data_in <= 24'b001001110011100101010000;
#10000;
data_in <= 24'b001010100011110001010011;
#10000;
data_in <= 24'b001001000011011101001100;
#10000;
data_in <= 24'b000110010010110001000001;
#10000;
data_in <= 24'b000100100010001100110110;
#10000;
data_in <= 24'b001000010011010001001111;
#10000;
data_in <= 24'b000111110011001001001101;
#10000;
data_in <= 24'b000111110011001001001101;
#10000;
data_in <= 24'b001001100011101001010011;
#10000;
data_in <= 24'b001011100100001001011011;
#10000;
data_in <= 24'b001100100100011101011101;
#10000;
data_in <= 24'b001011100100001101011001;
#10000;
data_in <= 24'b001010100011110101010010;
#10000;
data_in <= 24'b001001110011110001010111;
#10000;
data_in <= 24'b001000010011011001010001;
#10000;
data_in <= 24'b000111010011001001001101;
#10000;
data_in <= 24'b001000110011100001010011;
#10000;
data_in <= 24'b001100010100011101100000;
#10000;
data_in <= 24'b001111100101010001101101;
#10000;
data_in <= 24'b010000100101100101101111;
#10000;
data_in <= 24'b010001000101100101101111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001000110011001101000100;
#10000;
data_in <= 24'b001001110011100001001011;
#10000;
data_in <= 24'b001000010011001001000101;
#10000;
data_in <= 24'b000110000010101101000000;
#10000;
data_in <= 24'b001000110011011001001011;
#10000;
data_in <= 24'b001011110100001001010111;
#10000;
data_in <= 24'b001100110100010101011100;
#10000;
data_in <= 24'b001101100100100101011110;
#10000;
data_in <= 24'b000111000010101000111100;
#10000;
data_in <= 24'b000111100010111101000010;
#10000;
data_in <= 24'b000100110010010000110111;
#10000;
data_in <= 24'b000010010001101000101101;
#10000;
data_in <= 24'b000110010010101000111111;
#10000;
data_in <= 24'b001010010011110001010001;
#10000;
data_in <= 24'b001011000011111101010100;
#10000;
data_in <= 24'b001010000011101101010000;
#10000;
data_in <= 24'b000101100010010000110110;
#10000;
data_in <= 24'b000110010010100000111011;
#10000;
data_in <= 24'b000011010001110000101111;
#10000;
data_in <= 24'b000000110001010000100111;
#10000;
data_in <= 24'b000101000010010100111010;
#10000;
data_in <= 24'b001001110011100001001101;
#10000;
data_in <= 24'b001001100011011101001010;
#10000;
data_in <= 24'b001000000011000101000100;
#10000;
data_in <= 24'b000011110001110100110000;
#10000;
data_in <= 24'b000101000010001100110110;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b000110010010101000111111;
#10000;
data_in <= 24'b000111000010110101000010;
#10000;
data_in <= 24'b000110100010101100111110;
#10000;
data_in <= 24'b000110110010110000111111;
#10000;
data_in <= 24'b000010010001011100101010;
#10000;
data_in <= 24'b000100010001111100110010;
#10000;
data_in <= 24'b000110010010011100111101;
#10000;
data_in <= 24'b001000000010111001000100;
#10000;
data_in <= 24'b000111100010110001000010;
#10000;
data_in <= 24'b000011110001110100110011;
#10000;
data_in <= 24'b000010110001101000101101;
#10000;
data_in <= 24'b000110010010100000111011;
#10000;
data_in <= 24'b000101010010010000110111;
#10000;
data_in <= 24'b000111100010110000111111;
#10000;
data_in <= 24'b001000110011000101000111;
#10000;
data_in <= 24'b001001100011010001001010;
#10000;
data_in <= 24'b000111100010110001000010;
#10000;
data_in <= 24'b000010100001100000101110;
#10000;
data_in <= 24'b000010000001011100101010;
#10000;
data_in <= 24'b000110100010101000111011;
#10000;
data_in <= 24'b001100010011111101010101;
#10000;
data_in <= 24'b001101010100001001011000;
#10000;
data_in <= 24'b001010100011100001001110;
#10000;
data_in <= 24'b000111010010101101000001;
#10000;
data_in <= 24'b000110000010011000111100;
#10000;
data_in <= 24'b000100110010000100110111;
#10000;
data_in <= 24'b000100110010001000110101;
#10000;
data_in <= 24'b000111000010110000111101;
#10000;
data_in <= 24'b010001010101001101101001;
#10000;
data_in <= 24'b010001000101000101100111;
#10000;
data_in <= 24'b001010010011011101001101;
#10000;
data_in <= 24'b000011100001110000110010;
#10000;
data_in <= 24'b000011100001110000110010;
#10000;
data_in <= 24'b000110100010100000111110;
#10000;
data_in <= 24'b000111000010101100111110;
#10000;
data_in <= 24'b000110100010101000111011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001101100100100001011111;
#10000;
data_in <= 24'b001011000011111101010100;
#10000;
data_in <= 24'b000110110010110000111111;
#10000;
data_in <= 24'b000010010001100100101010;
#10000;
data_in <= 24'b000000000000111000011110;
#10000;
data_in <= 24'b000000000000101100011011;
#10000;
data_in <= 24'b000000000000100100010111;
#10000;
data_in <= 24'b000000000000010100010101;
#10000;
data_in <= 24'b001101000100011101011100;
#10000;
data_in <= 24'b001011110100000001010011;
#10000;
data_in <= 24'b001000000011000001000001;
#10000;
data_in <= 24'b000011010001110000101100;
#10000;
data_in <= 24'b000000100000111100011101;
#10000;
data_in <= 24'b000000000000101100010111;
#10000;
data_in <= 24'b000000000000100100010101;
#10000;
data_in <= 24'b000000000000011100010011;
#10000;
data_in <= 24'b001100000100000101010100;
#10000;
data_in <= 24'b001011110011111101010000;
#10000;
data_in <= 24'b001001000011010001000100;
#10000;
data_in <= 24'b000100100010001000101111;
#10000;
data_in <= 24'b000001000001001100011100;
#10000;
data_in <= 24'b000000000000110000010100;
#10000;
data_in <= 24'b000000000000101000010010;
#10000;
data_in <= 24'b000000000000101000010010;
#10000;
data_in <= 24'b001001100011011001000111;
#10000;
data_in <= 24'b001010010011100001001000;
#10000;
data_in <= 24'b001001000011010001000001;
#10000;
data_in <= 24'b000101110010010100110001;
#10000;
data_in <= 24'b000010010001010100011111;
#10000;
data_in <= 24'b000000110000111100010101;
#10000;
data_in <= 24'b000000010000101100010010;
#10000;
data_in <= 24'b000000000000101000010001;
#10000;
data_in <= 24'b000111000010101000111100;
#10000;
data_in <= 24'b000111110010111000111110;
#10000;
data_in <= 24'b000111100010101100111001;
#10000;
data_in <= 24'b000101100010001000101100;
#10000;
data_in <= 24'b000011010001100000100000;
#10000;
data_in <= 24'b000010000001001000011001;
#10000;
data_in <= 24'b000000110000110100010100;
#10000;
data_in <= 24'b000000100000101100001111;
#10000;
data_in <= 24'b000110000010011000111000;
#10000;
data_in <= 24'b000101110010011100110100;
#10000;
data_in <= 24'b000101100010001000101110;
#10000;
data_in <= 24'b000100010001101100100101;
#10000;
data_in <= 24'b000011100001011100100000;
#10000;
data_in <= 24'b000011000001011000011101;
#10000;
data_in <= 24'b000010010001001000010110;
#10000;
data_in <= 24'b000001000000110100010000;
#10000;
data_in <= 24'b000111010010101100111101;
#10000;
data_in <= 24'b000101000010010000110001;
#10000;
data_in <= 24'b000010110001011100100011;
#10000;
data_in <= 24'b000001100001000000011010;
#10000;
data_in <= 24'b000010100001001100011100;
#10000;
data_in <= 24'b000100010001100100100000;
#10000;
data_in <= 24'b000100000001011000011011;
#10000;
data_in <= 24'b000010010001000000010011;
#10000;
data_in <= 24'b001001000011001001000100;
#10000;
data_in <= 24'b000101000010010000110001;
#10000;
data_in <= 24'b000001010001000100011101;
#10000;
data_in <= 24'b000000000000101000010010;
#10000;
data_in <= 24'b000001110001000000011001;
#10000;
data_in <= 24'b000100110001110000100000;
#10000;
data_in <= 24'b000100110001100100011110;
#10000;
data_in <= 24'b000011000001010000010100;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000101100010001100111001;
#10000;
data_in <= 24'b001100110100000101011000;
#10000;
data_in <= 24'b010100100110000101111011;
#10000;
data_in <= 24'b010111010110111010001000;
#10000;
data_in <= 24'b010101110110100010000011;
#10000;
data_in <= 24'b010100010110011010000010;
#10000;
data_in <= 24'b010111100111001010010001;
#10000;
data_in <= 24'b011010101000000010100011;
#10000;
data_in <= 24'b000000000000011000010110;
#10000;
data_in <= 24'b000011010001101100101110;
#10000;
data_in <= 24'b001011010011101101001110;
#10000;
data_in <= 24'b010010100101100001101110;
#10000;
data_in <= 24'b010110010110101001111111;
#10000;
data_in <= 24'b010111000110111010000101;
#10000;
data_in <= 24'b010110010110101010000101;
#10000;
data_in <= 24'b010100010110011010000010;
#10000;
data_in <= 24'b000000000000000100001110;
#10000;
data_in <= 24'b000000000000010100010011;
#10000;
data_in <= 24'b000010000001001100100001;
#10000;
data_in <= 24'b000111110010110000111100;
#10000;
data_in <= 24'b001110010100011101011001;
#10000;
data_in <= 24'b010011010101110001101111;
#10000;
data_in <= 24'b010101000110001001111001;
#10000;
data_in <= 24'b010011110110000001111010;
#10000;
data_in <= 24'b000000000000100100010010;
#10000;
data_in <= 24'b000000000000100000010000;
#10000;
data_in <= 24'b000000000000010100001111;
#10000;
data_in <= 24'b000000000000100100010011;
#10000;
data_in <= 24'b000011000001011100100101;
#10000;
data_in <= 24'b001000010010111000111110;
#10000;
data_in <= 24'b001110000100011001011000;
#10000;
data_in <= 24'b010010000101011101101010;
#10000;
data_in <= 24'b000000000000010000001000;
#10000;
data_in <= 24'b000000000000100000001100;
#10000;
data_in <= 24'b000000000000100000001111;
#10000;
data_in <= 24'b000000000000011000001101;
#10000;
data_in <= 24'b000000000000001100001101;
#10000;
data_in <= 24'b000000010000101000010111;
#10000;
data_in <= 24'b000011110001101000101000;
#10000;
data_in <= 24'b000110100010011100110111;
#10000;
data_in <= 24'b000000010000100000001011;
#10000;
data_in <= 24'b000000100000100100001100;
#10000;
data_in <= 24'b000000110000101000001101;
#10000;
data_in <= 24'b000000000000100100001101;
#10000;
data_in <= 24'b000000000000011000001101;
#10000;
data_in <= 24'b000000000000010000001101;
#10000;
data_in <= 24'b000000000000001100001101;
#10000;
data_in <= 24'b000000000000001100001111;
#10000;
data_in <= 24'b000011110001010000010101;
#10000;
data_in <= 24'b000010000001000000010000;
#10000;
data_in <= 24'b000000110000101100001011;
#10000;
data_in <= 24'b000000000000100100001001;
#10000;
data_in <= 24'b000000000000100100001100;
#10000;
data_in <= 24'b000000000000100100001101;
#10000;
data_in <= 24'b000000000000011000001101;
#10000;
data_in <= 24'b000000000000001100001011;
#10000;
data_in <= 24'b000011010001001000010011;
#10000;
data_in <= 24'b000010110001000100010000;
#10000;
data_in <= 24'b000001100000111000001101;
#10000;
data_in <= 24'b000001000000110000001011;
#10000;
data_in <= 24'b000000010000101000001101;
#10000;
data_in <= 24'b000000000000100100001100;
#10000;
data_in <= 24'b000000000000100000001111;
#10000;
data_in <= 24'b000000000000100000001111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011001110111111110100011;
#10000;
data_in <= 24'b011000100111110010100001;
#10000;
data_in <= 24'b011000010111101110100011;
#10000;
data_in <= 24'b011000010111110110100110;
#10000;
data_in <= 24'b011000100111111110101011;
#10000;
data_in <= 24'b011000101000000110101110;
#10000;
data_in <= 24'b011001001000001110110000;
#10000;
data_in <= 24'b011001111000011110110010;
#10000;
data_in <= 24'b010101000110100110001001;
#10000;
data_in <= 24'b010101010110111010010000;
#10000;
data_in <= 24'b010111010111010110011001;
#10000;
data_in <= 24'b011000010111101110100000;
#10000;
data_in <= 24'b011001101000000010101000;
#10000;
data_in <= 24'b011001101000001010101011;
#10000;
data_in <= 24'b011001011000000010101100;
#10000;
data_in <= 24'b011000010111111110101000;
#10000;
data_in <= 24'b010011010101111101111100;
#10000;
data_in <= 24'b010100010110011010000101;
#10000;
data_in <= 24'b010101010110101010001010;
#10000;
data_in <= 24'b010100110110100110001100;
#10000;
data_in <= 24'b010101010110110110010001;
#10000;
data_in <= 24'b010111000111011010011010;
#10000;
data_in <= 24'b011000100111110010100001;
#10000;
data_in <= 24'b011000000111101110100000;
#10000;
data_in <= 24'b010010010101100101110000;
#10000;
data_in <= 24'b010011110110000001111010;
#10000;
data_in <= 24'b010100000110001101111110;
#10000;
data_in <= 24'b010010010101111001111010;
#10000;
data_in <= 24'b010010110101111101111110;
#10000;
data_in <= 24'b010101010110101010001010;
#10000;
data_in <= 24'b010111010111001010010010;
#10000;
data_in <= 24'b010110010111001010010100;
#10000;
data_in <= 24'b001001110011010101000111;
#10000;
data_in <= 24'b001101010100010001010111;
#10000;
data_in <= 24'b010000000101000101100110;
#10000;
data_in <= 24'b010000110101010101101100;
#10000;
data_in <= 24'b010001110101100001110010;
#10000;
data_in <= 24'b010011000101111101111010;
#10000;
data_in <= 24'b010100000110001101111110;
#10000;
data_in <= 24'b010011010110001010000001;
#10000;
data_in <= 24'b000000100000111100011101;
#10000;
data_in <= 24'b000010100001100100101001;
#10000;
data_in <= 24'b000101110010010100110111;
#10000;
data_in <= 24'b000111110010111001000001;
#10000;
data_in <= 24'b001001100011010001001010;
#10000;
data_in <= 24'b001011110100000001010101;
#10000;
data_in <= 24'b001111100100111001100101;
#10000;
data_in <= 24'b010001010101100001110011;
#10000;
data_in <= 24'b000000000000010100001111;
#10000;
data_in <= 24'b000000000000001100001111;
#10000;
data_in <= 24'b000000000000010000010010;
#10000;
data_in <= 24'b000000000000100100011001;
#10000;
data_in <= 24'b000000010000110100011111;
#10000;
data_in <= 24'b000010010001011100101001;
#10000;
data_in <= 24'b001000010010111101000010;
#10000;
data_in <= 24'b001101100100011001011101;
#10000;
data_in <= 24'b000000000000101000010100;
#10000;
data_in <= 24'b000000000000010000001110;
#10000;
data_in <= 24'b000000000000001100010001;
#10000;
data_in <= 24'b000000000000100000010110;
#10000;
data_in <= 24'b000000000000010100010101;
#10000;
data_in <= 24'b000000000000010100010101;
#10000;
data_in <= 24'b000010000001011000101000;
#10000;
data_in <= 24'b000111010010111001000011;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b011011001000110110110100;
#10000;
data_in <= 24'b011011001001000010110100;
#10000;
data_in <= 24'b011011011001000110110111;
#10000;
data_in <= 24'b011011101001001110111001;
#10000;
data_in <= 24'b011100011001010110111101;
#10000;
data_in <= 24'b011101001001101111000010;
#10000;
data_in <= 24'b011110001010000011001010;
#10000;
data_in <= 24'b011111001010010011001110;
#10000;
data_in <= 24'b011010001000011110101110;
#10000;
data_in <= 24'b011010001000101010101110;
#10000;
data_in <= 24'b011010101000101110110010;
#10000;
data_in <= 24'b011010101000111010110100;
#10000;
data_in <= 24'b011011011001000010111000;
#10000;
data_in <= 24'b011100001001010010111100;
#10000;
data_in <= 24'b011100111001100111000011;
#10000;
data_in <= 24'b011101011001110111000111;
#10000;
data_in <= 24'b011000100111111110100100;
#10000;
data_in <= 24'b011000111000001110100110;
#10000;
data_in <= 24'b011001101000011010101010;
#10000;
data_in <= 24'b011001111000100110101101;
#10000;
data_in <= 24'b011010001000110010110010;
#10000;
data_in <= 24'b011010101000111110110101;
#10000;
data_in <= 24'b011011101001001010111010;
#10000;
data_in <= 24'b011011101001010110111100;
#10000;
data_in <= 24'b010110100111011010011001;
#10000;
data_in <= 24'b010110110111100110011100;
#10000;
data_in <= 24'b011000000111110110100010;
#10000;
data_in <= 24'b011000101000001010100110;
#10000;
data_in <= 24'b011000111000010010101011;
#10000;
data_in <= 24'b011001001000100010101110;
#10000;
data_in <= 24'b011001111000101010110010;
#10000;
data_in <= 24'b011010001000110010110100;
#10000;
data_in <= 24'b010011100110011110001001;
#10000;
data_in <= 24'b010011110110101110001110;
#10000;
data_in <= 24'b010101010111000110010100;
#10000;
data_in <= 24'b010101110111010110011000;
#10000;
data_in <= 24'b010110010111100110011101;
#10000;
data_in <= 24'b010110100111110010100000;
#10000;
data_in <= 24'b010111010111111010100101;
#10000;
data_in <= 24'b010111011000000110100111;
#10000;
data_in <= 24'b001111110101011001110110;
#10000;
data_in <= 24'b001111100101100001111100;
#10000;
data_in <= 24'b010000110101110110000001;
#10000;
data_in <= 24'b010001100110001010000101;
#10000;
data_in <= 24'b010001110110010010001001;
#10000;
data_in <= 24'b010010000110100010001100;
#10000;
data_in <= 24'b010010100110100110010000;
#10000;
data_in <= 24'b010010100110101110010010;
#10000;
data_in <= 24'b001100110100100001101000;
#10000;
data_in <= 24'b001100100100101001101110;
#10000;
data_in <= 24'b001101010100110101110001;
#10000;
data_in <= 24'b001101010100111101110011;
#10000;
data_in <= 24'b001101010101000101110100;
#10000;
data_in <= 24'b001101010101001101110110;
#10000;
data_in <= 24'b001101010101010101111001;
#10000;
data_in <= 24'b001101010101011001111101;
#10000;
data_in <= 24'b001011100100000101100010;
#10000;
data_in <= 24'b001011000100001001100110;
#10000;
data_in <= 24'b001011000100010001101000;
#10000;
data_in <= 24'b001010110100010101101001;
#10000;
data_in <= 24'b001010110100010101101001;
#10000;
data_in <= 24'b001010000100011001101001;
#10000;
data_in <= 24'b001010100100011101101100;
#10000;
data_in <= 24'b001010010100100101101101;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100001001010110011010110;
#10000;
data_in <= 24'b100010001011000011011010;
#10000;
data_in <= 24'b100011101011010011011110;
#10000;
data_in <= 24'b100100001011011111011110;
#10000;
data_in <= 24'b100101101011101011100010;
#10000;
data_in <= 24'b100110101011111111100101;
#10000;
data_in <= 24'b100110101011111011100100;
#10000;
data_in <= 24'b100101101011101011100000;
#10000;
data_in <= 24'b011110111010000111001011;
#10000;
data_in <= 24'b100000001010011011010000;
#10000;
data_in <= 24'b100001001010101011010100;
#10000;
data_in <= 24'b100001101010110011010110;
#10000;
data_in <= 24'b100010111010111111010111;
#10000;
data_in <= 24'b100011011011000111011001;
#10000;
data_in <= 24'b100011001010111111010111;
#10000;
data_in <= 24'b100001101010100111010001;
#10000;
data_in <= 24'b011100111001011011000001;
#10000;
data_in <= 24'b011110001001101111000110;
#10000;
data_in <= 24'b011111001001111111001010;
#10000;
data_in <= 24'b011111101010000111001100;
#10000;
data_in <= 24'b100000001010001011001101;
#10000;
data_in <= 24'b011111111010000111001100;
#10000;
data_in <= 24'b011110111001101111000110;
#10000;
data_in <= 24'b011101001001010010111111;
#10000;
data_in <= 24'b011011001000111110111010;
#10000;
data_in <= 24'b011100011001010010111111;
#10000;
data_in <= 24'b011101011001100011000011;
#10000;
data_in <= 24'b011101011001100011000011;
#10000;
data_in <= 24'b011101011001011111000010;
#10000;
data_in <= 24'b011100011001001010111111;
#10000;
data_in <= 24'b011010101000100110110110;
#10000;
data_in <= 24'b011000011000000010101101;
#10000;
data_in <= 24'b011000011000010010101100;
#10000;
data_in <= 24'b011001011000100010110000;
#10000;
data_in <= 24'b011010001000101010110101;
#10000;
data_in <= 24'b011001111000100110110100;
#10000;
data_in <= 24'b011001011000010010110001;
#10000;
data_in <= 24'b011000000111111010101101;
#10000;
data_in <= 24'b010110000111010010100011;
#10000;
data_in <= 24'b010011100110101110011000;
#10000;
data_in <= 24'b010011010110110110010110;
#10000;
data_in <= 24'b010011110111001010011010;
#10000;
data_in <= 24'b010100000111001010011101;
#10000;
data_in <= 24'b010011100110111110011100;
#10000;
data_in <= 24'b010011010110101110011010;
#10000;
data_in <= 24'b010010010110011110010110;
#10000;
data_in <= 24'b010000100101111010001101;
#10000;
data_in <= 24'b001110010101010110000100;
#10000;
data_in <= 24'b001101110101011110000000;
#10000;
data_in <= 24'b001110100101101010000011;
#10000;
data_in <= 24'b001110110101101110000110;
#10000;
data_in <= 24'b001110010101100010000101;
#10000;
data_in <= 24'b001110100101011010000101;
#10000;
data_in <= 24'b001110000101010010000011;
#10000;
data_in <= 24'b001101000100110101111111;
#10000;
data_in <= 24'b001011010100011101110110;
#10000;
data_in <= 24'b001010110100101101110100;
#10000;
data_in <= 24'b001011010100110101110110;
#10000;
data_in <= 24'b001011100100110101111010;
#10000;
data_in <= 24'b001011010100110001111001;
#10000;
data_in <= 24'b001100000100110001111011;
#10000;
data_in <= 24'b001100000100110001111011;
#10000;
data_in <= 24'b001011110100100001111010;
#10000;
data_in <= 24'b001010010100001101110010;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b100011001011000011010110;
#10000;
data_in <= 24'b100010011010110011010100;
#10000;
data_in <= 24'b100000101010010111001101;
#10000;
data_in <= 24'b011110011001101111000110;
#10000;
data_in <= 24'b011011001000110110111010;
#10000;
data_in <= 24'b010110010111101010100111;
#10000;
data_in <= 24'b010010000110011010010101;
#10000;
data_in <= 24'b001110110101100110001000;
#10000;
data_in <= 24'b100001011010100011010000;
#10000;
data_in <= 24'b011111011010000011001000;
#10000;
data_in <= 24'b011011101001000010111011;
#10000;
data_in <= 24'b010111111000000110101100;
#10000;
data_in <= 24'b010011110111000010011101;
#10000;
data_in <= 24'b010000010110000010001101;
#10000;
data_in <= 24'b001100100101000001111111;
#10000;
data_in <= 24'b001010100100011101110100;
#10000;
data_in <= 24'b011100001001001010111101;
#10000;
data_in <= 24'b011000111000010110110000;
#10000;
data_in <= 24'b010100100111000110011110;
#10000;
data_in <= 24'b001111110101111010001011;
#10000;
data_in <= 24'b001100010101000001111101;
#10000;
data_in <= 24'b001010010100011001110011;
#10000;
data_in <= 24'b001000010011111001101011;
#10000;
data_in <= 24'b000111110011100101100111;
#10000;
data_in <= 24'b010100110111001110011110;
#10000;
data_in <= 24'b010010000110100010010011;
#10000;
data_in <= 24'b001101110101011010000011;
#10000;
data_in <= 24'b001010010100100001110101;
#10000;
data_in <= 24'b001000110100000001101101;
#10000;
data_in <= 24'b001000100011110001101010;
#10000;
data_in <= 24'b001000010011101101101001;
#10000;
data_in <= 24'b001000100011101101100111;
#10000;
data_in <= 24'b001111010101101010000110;
#10000;
data_in <= 24'b001101010101001001111110;
#10000;
data_in <= 24'b001011000100100101110101;
#10000;
data_in <= 24'b001001000100000101101101;
#10000;
data_in <= 24'b001000110011111001101010;
#10000;
data_in <= 24'b001000100011110101101001;
#10000;
data_in <= 24'b001000100011101101100111;
#10000;
data_in <= 24'b001000100011100101100110;
#10000;
data_in <= 24'b001100010100111001111011;
#10000;
data_in <= 24'b001011000100100101110101;
#10000;
data_in <= 24'b001001110100010001110000;
#10000;
data_in <= 24'b001001010100000001101100;
#10000;
data_in <= 24'b001000100011110101101001;
#10000;
data_in <= 24'b001000010011101001100110;
#10000;
data_in <= 24'b000111100011010101100010;
#10000;
data_in <= 24'b000110100011001001011100;
#10000;
data_in <= 24'b001011000100011001110100;
#10000;
data_in <= 24'b001010010100010001110000;
#10000;
data_in <= 24'b001001000011111101101011;
#10000;
data_in <= 24'b001000010011110001101000;
#10000;
data_in <= 24'b001000100011101101100111;
#10000;
data_in <= 24'b001000000011011101100100;
#10000;
data_in <= 24'b000111000011010001011110;
#10000;
data_in <= 24'b000110100011000001011010;
#10000;
data_in <= 24'b001001110100000101101111;
#10000;
data_in <= 24'b001000110011111001101010;
#10000;
data_in <= 24'b000111110011101001100110;
#10000;
data_in <= 24'b000111010011100001100100;
#10000;
data_in <= 24'b001000000011011101100100;
#10000;
data_in <= 24'b001000010011100001100101;
#10000;
data_in <= 24'b001000010011011101100001;
#10000;
data_in <= 24'b000111110011010101011111;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b001011010100101001110111;
#10000;
data_in <= 24'b001010100100011001101111;
#10000;
data_in <= 24'b001001100011111101100111;
#10000;
data_in <= 24'b000111110011011101011011;
#10000;
data_in <= 24'b000110100011000101010001;
#10000;
data_in <= 24'b000101000010100101001000;
#10000;
data_in <= 24'b000011110010010001000000;
#10000;
data_in <= 24'b000011110010000000111010;
#10000;
data_in <= 24'b001010010100010001110000;
#10000;
data_in <= 24'b001001110100000001101010;
#10000;
data_in <= 24'b001000110011100101100010;
#10000;
data_in <= 24'b000111010011001101010111;
#10000;
data_in <= 24'b000110010010111001001110;
#10000;
data_in <= 24'b000100100010011101000110;
#10000;
data_in <= 24'b000011010010001000111110;
#10000;
data_in <= 24'b000011010001111000111000;
#10000;
data_in <= 24'b001000110011110001101000;
#10000;
data_in <= 24'b001000000011100101100001;
#10000;
data_in <= 24'b000111000011001101011001;
#10000;
data_in <= 24'b000110000010111001010001;
#10000;
data_in <= 24'b000101010010101001001010;
#10000;
data_in <= 24'b000100000010010101000100;
#10000;
data_in <= 24'b000011000010000100111101;
#10000;
data_in <= 24'b000010110001111000111001;
#10000;
data_in <= 24'b000111010011010101011111;
#10000;
data_in <= 24'b000111000011001001011011;
#10000;
data_in <= 24'b000110010010111001010100;
#10000;
data_in <= 24'b000101010010101101001110;
#10000;
data_in <= 24'b000101000010100101001001;
#10000;
data_in <= 24'b000100000010010101000100;
#10000;
data_in <= 24'b000011100010001001000001;
#10000;
data_in <= 24'b000010110010000000111011;
#10000;
data_in <= 24'b000110100011001001011100;
#10000;
data_in <= 24'b000110010010111101011000;
#10000;
data_in <= 24'b000110000010110101010011;
#10000;
data_in <= 24'b000101010010101101001110;
#10000;
data_in <= 24'b000101100010101101001011;
#10000;
data_in <= 24'b000101000010100101001000;
#10000;
data_in <= 24'b000100010010011001000101;
#10000;
data_in <= 24'b000100010010011001000010;
#10000;
data_in <= 24'b000110110011000101011011;
#10000;
data_in <= 24'b000110010010111101011000;
#10000;
data_in <= 24'b000110000010110101010011;
#10000;
data_in <= 24'b000101110010110101010001;
#10000;
data_in <= 24'b000110010010110101010000;
#10000;
data_in <= 24'b000110000010110101001101;
#10000;
data_in <= 24'b000101110010110001001100;
#10000;
data_in <= 24'b000101010010101101000111;
#10000;
data_in <= 24'b000110110011000101011011;
#10000;
data_in <= 24'b000110010010111101011000;
#10000;
data_in <= 24'b000110010010111001010100;
#10000;
data_in <= 24'b000110010010111101010011;
#10000;
data_in <= 24'b000110010010111101010010;
#10000;
data_in <= 24'b000110010011000001010000;
#10000;
data_in <= 24'b000110010011000001010000;
#10000;
data_in <= 24'b000110100010111101001110;
#10000;
data_in <= 24'b000110110011000101011010;
#10000;
data_in <= 24'b000110010010111101011000;
#10000;
data_in <= 24'b000110100010111101010101;
#10000;
data_in <= 24'b000110100011000001010100;
#10000;
data_in <= 24'b000110100011000001010100;
#10000;
data_in <= 24'b000110110011000101010100;
#10000;
data_in <= 24'b000110110011001001010010;
#10000;
data_in <= 24'b000110100011001001010000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
data_in <= 24'b000100000001111000110101;
#10000;
data_in <= 24'b000100010001111000110100;
#10000;
data_in <= 24'b000100000001111000110001;
#10000;
data_in <= 24'b000100000001111000110000;
#10000;
data_in <= 24'b000100110001111100110001;
#10000;
data_in <= 24'b000100110010000000101110;
#10000;
data_in <= 24'b000101100010000100101111;
#10000;
data_in <= 24'b000101110010001100101111;
#10000;
data_in <= 24'b000100000001111000110101;
#10000;
data_in <= 24'b000100010001111000110100;
#10000;
data_in <= 24'b000100010001111100110010;
#10000;
data_in <= 24'b000100010001111100110010;
#10000;
data_in <= 24'b000100110001111100110001;
#10000;
data_in <= 24'b000101000010000100110001;
#10000;
data_in <= 24'b000101110010001000110000;
#10000;
data_in <= 24'b000101110010001100101111;
#10000;
data_in <= 24'b000100000001111100111001;
#10000;
data_in <= 24'b000100100010000000110110;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b000100100010000000110010;
#10000;
data_in <= 24'b000100110010001000110010;
#10000;
data_in <= 24'b000101010010001000110000;
#10000;
data_in <= 24'b000101100010001100110001;
#10000;
data_in <= 24'b000100010010001000111100;
#10000;
data_in <= 24'b000100110010001100111010;
#10000;
data_in <= 24'b000100100010001100111000;
#10000;
data_in <= 24'b000100110010001000110101;
#10000;
data_in <= 24'b000100110010001000110101;
#10000;
data_in <= 24'b000101000010001000110100;
#10000;
data_in <= 24'b000101100010001100110011;
#10000;
data_in <= 24'b000101110010010000110010;
#10000;
data_in <= 24'b000101000010011101000010;
#10000;
data_in <= 24'b000101010010011100111110;
#10000;
data_in <= 24'b000101000010011000111101;
#10000;
data_in <= 24'b000101000010010100111010;
#10000;
data_in <= 24'b000101010010010000110111;
#10000;
data_in <= 24'b000101100010010000110110;
#10000;
data_in <= 24'b000101110010001100110101;
#10000;
data_in <= 24'b000101110010010000110100;
#10000;
data_in <= 24'b000101110010110001000111;
#10000;
data_in <= 24'b000110000010110001000101;
#10000;
data_in <= 24'b000101100010101001000011;
#10000;
data_in <= 24'b000101100010100000111111;
#10000;
data_in <= 24'b000101100010011100111100;
#10000;
data_in <= 24'b000101100010010100111000;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
data_in <= 24'b000110000010010000110110;
#10000;
data_in <= 24'b000110110011000101001101;
#10000;
data_in <= 24'b000110110011000101001010;
#10000;
data_in <= 24'b000110100010111001000111;
#10000;
data_in <= 24'b000110010010101101000010;
#10000;
data_in <= 24'b000110000010100100111110;
#10000;
data_in <= 24'b000110000010011100111010;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
data_in <= 24'b000111100011010001010000;
#10000;
data_in <= 24'b000111010011010001001110;
#10000;
data_in <= 24'b000111010011000101001010;
#10000;
data_in <= 24'b000110010010111001000100;
#10000;
data_in <= 24'b000110100010101001000001;
#10000;
data_in <= 24'b000101110010100000111101;
#10000;
data_in <= 24'b000110000010011000111001;
#10000;
data_in <= 24'b000101110010010100111000;
#10000;
#130000;
enable <= 1'b0;
#10000;
enable <= 1'b1;
end_of_file_signal  <= 1'b1;
data_in <= 24'b000101100010001000101100;
#10000;
data_in <= 24'b000110000010010000101110;
#10000;
data_in <= 24'b000101100010010100101110;
#10000;
data_in <= 24'b000100100010001100101100;
#10000;
data_in <= 24'b000011110010000100101100;
#10000;
data_in <= 24'b000100000010001000101101;
#10000;
data_in <= 24'b000100000010001100110000;
#10000;
data_in <= 24'b000011110010010100110001;
#10000;
data_in <= 24'b000101110010001100101111;
#10000;
data_in <= 24'b000101010010010000101101;
#10000;
data_in <= 24'b000100110010000100101101;
#10000;
data_in <= 24'b000100000010000000101100;
#10000;
data_in <= 24'b000011100010000000101011;
#10000;
data_in <= 24'b000100000010000100101110;
#10000;
data_in <= 24'b000100010010010000110001;
#10000;
data_in <= 24'b000100000010011000110010;
#10000;
data_in <= 24'b000110010010011000110100;
#10000;
data_in <= 24'b000101010010001100101111;
#10000;
data_in <= 24'b000100100001111100101101;
#10000;
data_in <= 24'b000011110001111100101100;
#10000;
data_in <= 24'b000100000010000100101110;
#10000;
data_in <= 24'b000100100010001000110010;
#10000;
data_in <= 24'b000100100010010100110100;
#10000;
data_in <= 24'b000100110010011000110101;
#10000;
data_in <= 24'b000110100010011100110111;
#10000;
data_in <= 24'b000101100010001100110001;
#10000;
data_in <= 24'b000100100001111100101111;
#10000;
data_in <= 24'b000100110010000000110000;
#10000;
data_in <= 24'b000100110010001000110010;
#10000;
data_in <= 24'b000100100010001000110011;
#10000;
data_in <= 24'b000100110010001100110100;
#10000;
data_in <= 24'b000100100010010000110101;
#10000;
data_in <= 24'b000110000010010000110110;
#10000;
data_in <= 24'b000101000010000100110001;
#10000;
data_in <= 24'b000100100001111000110000;
#10000;
data_in <= 24'b000101010010000100110011;
#10000;
data_in <= 24'b000101100010001000110100;
#10000;
data_in <= 24'b000100010001111100110010;
#10000;
data_in <= 24'b000100000001111000110001;
#10000;
data_in <= 24'b000100010010000000110011;
#10000;
data_in <= 24'b000101100010001000110100;
#10000;
data_in <= 24'b000100100001111000110000;
#10000;
data_in <= 24'b000100100001111000110000;
#10000;
data_in <= 24'b000101100010000100110101;
#10000;
data_in <= 24'b000101000001111100110011;
#10000;
data_in <= 24'b000100000001101100110001;
#10000;
data_in <= 24'b000100000001110100110011;
#10000;
data_in <= 24'b000101100010001100111001;
#10000;
data_in <= 24'b000101110010001000110110;
#10000;
data_in <= 24'b000101000001111100110011;
#10000;
data_in <= 24'b000101110010000000110100;
#10000;
data_in <= 24'b000110100010001100110111;
#10000;
data_in <= 24'b000101010010000000110110;
#10000;
data_in <= 24'b000100100001110000110100;
#10000;
data_in <= 24'b000110010010001100111011;
#10000;
data_in <= 24'b001001010010111101000111;
#10000;
data_in <= 24'b000110110010011000111010;
#10000;
data_in <= 24'b000110000010001100110111;
#10000;
data_in <= 24'b000110100010001100110111;
#10000;
data_in <= 24'b000111010010011000111010;
#10000;
data_in <= 24'b000110000010001000111010;
#10000;
data_in <= 24'b000101100010000000111000;
#10000;
data_in <= 24'b001000100010101101000110;
#10000;
data_in <= 24'b001100110011110001010111;
#10000;
#130000;
enable <= 1'b0;

#2000000; 

$finish;
end // end of stimulus process
	
always
begin : CLOCK_clk
	//this process was generated based on formula: 0 0 ns, 1 5 ns -r 10 ns
	//#<time to next event>; // <current time>
	clk = 1'b0;
	#5000; //0
	clk = 1'b1;
	#5000; //5000
end

always 	@(JPEG_bitstream or data_ready)
begin : JPEG
		if (data_ready==1'b1) 		
					$display("%h", JPEG_bitstream);						
end	


endmodule
